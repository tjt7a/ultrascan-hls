




/*
******************** Summary ********************
report for vasim_50
Number of nodes = 258
Number of edges = 258
Average edge per node = 1.0
Number of start nodes = 1
Number of report nodes = 1
does have all_input = True
does have special element = False
is Homogenous = True
stride value = 1
Max Fan-in = 2
Max Fan-out = 2
Max value in dim = 255
average number of intervals per STE = 1.96899224806
#######################################################
*/

 



module LUT_Match_vasim_50_1 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_2 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_3 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_4 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_5 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_6 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_7 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_8 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_9 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_10 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_11 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_12 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_13 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_14 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_15 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_16 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_17 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_18 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_19 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_20 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_21 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_22 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_23 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_24 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_25 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_26 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_27 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_28 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_29 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_30 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_31 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_32 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_33 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_34 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_35 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_36 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_37 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_38 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_39 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_40 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_41 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_42 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_43 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_44 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_45 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_46 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_47 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_48 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_49 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_50 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_51 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_52 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_53 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_54 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_55 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_56 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_57 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_58 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_59 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_60 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_61 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_62 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_63 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_64 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_65 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_66 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_67 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_68 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_69 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_70 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_71 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_72 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_73 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_74 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_75 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_76 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_77 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_78 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_79 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_80 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_81 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_82 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_83 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_84 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_85 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_86 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_87 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_88 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_89 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_90 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_91 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_92 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_93 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_94 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_95 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_96 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_97 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_98 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_99 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_100 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_101 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_102 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_103 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_104 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_105 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_106 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_107 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_108 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_109 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_110 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_111 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_112 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_113 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_114 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_115 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_116 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_117 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_118 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_119 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_120 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_121 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_122 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_123 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_124 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_125 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_126 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_127 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_128 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_129 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_130 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_131 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_132 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_133 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_134 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_135 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_136 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_137 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_138 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_139 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_140 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_141 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_142 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_143 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_144 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_145 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_146 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_147 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_148 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_149 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_150 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_151 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_152 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_153 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_154 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_155 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_156 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_157 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_158 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_159 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_160 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_161 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_162 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_163 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_164 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_165 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_166 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_167 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_168 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_169 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_170 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_171 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_172 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_173 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_174 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_175 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd35) &&(input_capture[7:0] <= 8'd35) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_176 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd33) &&(input_capture[7:0] <= 8'd33) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_177 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_178 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd33) &&(input_capture[7:0] <= 8'd33) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_179 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd33) &&(input_capture[7:0] <= 8'd33) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_180 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_181 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_182 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_183 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_184 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_185 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_186 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_187 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_188 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_189 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_190 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_191 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_192 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_193 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd35) &&(input_capture[7:0] <= 8'd35) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_194 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_195 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_196 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_197 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_198 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_199 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_200 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_201 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_202 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_203 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_204 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd36) &&(input_capture[7:0] <= 8'd36) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_205 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_206 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_207 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_208 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_209 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_210 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_211 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_212 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_213 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_214 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_215 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd36) &&(input_capture[7:0] <= 8'd36) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_216 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_217 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_218 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_219 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_220 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_221 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_222 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_223 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_224 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_225 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_226 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd36) &&(input_capture[7:0] <= 8'd36) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_227 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_228 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_229 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_230 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_231 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_232 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_233 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_234 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_235 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_236 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_237 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_238 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_239 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_240 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_241 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_242 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_243 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_244 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_245 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_246 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_247 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_248 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_249 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_250 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_251 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_252 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_253 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_254 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_255 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_256 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_257 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule

 



module LUT_Match_vasim_50_258 #(parameter integer width = 8)(
        input clk,
        input [width-1:0] symbols,
        output match);

wire match_internal;
wire [width-1:0] input_capture;
assign input_capture = symbols;
assign match = match_internal;

assign match_internal = (((input_capture[7:0] >= 8'd48) &&(input_capture[7:0] <= 8'd57) && 1'b1) ||
     ((input_capture[7:0] >= 8'd65) &&(input_capture[7:0] <= 8'd70) && 1'b1) ||
      1'b0) ? 1'b1 : 1'b0;


endmodule



module Automata_vasim_50(input clk,
           input run,
           input reset,
           input [7 : 0] symbols
           
           , output vasim_50_w_out_179);

wire all_input;
wire start_of_data;

assign all_input = 1'b1;
assign start_of_data = ~reset;



/*wire vasim_50_w_out_1;
*/

wire vasim_50_lut_match_1;
wire vasim_50_w_match_1;

    
    
    

LUT_Match_vasim_50_1 #(8) lut_match_vasim_50_1(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_1));


assign vasim_50_w_match_1 = vasim_50_lut_match_1 ;

STE #(.fan_in(1)) vasim_50_ste_1 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_248 }),
                .match(vasim_50_w_match_1) ,
                .active_state(vasim_50_w_out_1));




/*wire vasim_50_w_out_2;
*/

wire vasim_50_lut_match_2;
wire vasim_50_w_match_2;

    
    
    

LUT_Match_vasim_50_2 #(8) lut_match_vasim_50_2(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_2));


assign vasim_50_w_match_2 = vasim_50_lut_match_2 ;

STE #(.fan_in(1)) vasim_50_ste_2 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_258 }),
                .match(vasim_50_w_match_2) ,
                .active_state(vasim_50_w_out_2));




/*wire vasim_50_w_out_3;
*/

wire vasim_50_lut_match_3;
wire vasim_50_w_match_3;

    
    
    

LUT_Match_vasim_50_3 #(8) lut_match_vasim_50_3(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_3));


assign vasim_50_w_match_3 = vasim_50_lut_match_3 ;

STE #(.fan_in(1)) vasim_50_ste_3 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_2 }),
                .match(vasim_50_w_match_3) ,
                .active_state(vasim_50_w_out_3));




/*wire vasim_50_w_out_4;
*/

wire vasim_50_lut_match_4;
wire vasim_50_w_match_4;

    
    
    

LUT_Match_vasim_50_4 #(8) lut_match_vasim_50_4(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_4));


assign vasim_50_w_match_4 = vasim_50_lut_match_4 ;

STE #(.fan_in(1)) vasim_50_ste_4 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_3 }),
                .match(vasim_50_w_match_4) ,
                .active_state(vasim_50_w_out_4));




/*wire vasim_50_w_out_5;
*/

wire vasim_50_lut_match_5;
wire vasim_50_w_match_5;

    
    
    

LUT_Match_vasim_50_5 #(8) lut_match_vasim_50_5(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_5));


assign vasim_50_w_match_5 = vasim_50_lut_match_5 ;

STE #(.fan_in(1)) vasim_50_ste_5 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_4 }),
                .match(vasim_50_w_match_5) ,
                .active_state(vasim_50_w_out_5));




/*wire vasim_50_w_out_6;
*/

wire vasim_50_lut_match_6;
wire vasim_50_w_match_6;

    
    
    

LUT_Match_vasim_50_6 #(8) lut_match_vasim_50_6(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_6));


assign vasim_50_w_match_6 = vasim_50_lut_match_6 ;

STE #(.fan_in(1)) vasim_50_ste_6 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_5 }),
                .match(vasim_50_w_match_6) ,
                .active_state(vasim_50_w_out_6));




/*wire vasim_50_w_out_7;
*/

wire vasim_50_lut_match_7;
wire vasim_50_w_match_7;

    
    
    

LUT_Match_vasim_50_7 #(8) lut_match_vasim_50_7(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_7));


assign vasim_50_w_match_7 = vasim_50_lut_match_7 ;

STE #(.fan_in(1)) vasim_50_ste_7 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_6 }),
                .match(vasim_50_w_match_7) ,
                .active_state(vasim_50_w_out_7));




/*wire vasim_50_w_out_8;
*/

wire vasim_50_lut_match_8;
wire vasim_50_w_match_8;

    
    
    

LUT_Match_vasim_50_8 #(8) lut_match_vasim_50_8(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_8));


assign vasim_50_w_match_8 = vasim_50_lut_match_8 ;

STE #(.fan_in(1)) vasim_50_ste_8 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_7 }),
                .match(vasim_50_w_match_8) ,
                .active_state(vasim_50_w_out_8));




/*wire vasim_50_w_out_9;
*/

wire vasim_50_lut_match_9;
wire vasim_50_w_match_9;

    
    
    

LUT_Match_vasim_50_9 #(8) lut_match_vasim_50_9(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_9));


assign vasim_50_w_match_9 = vasim_50_lut_match_9 ;

STE #(.fan_in(1)) vasim_50_ste_9 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_8 }),
                .match(vasim_50_w_match_9) ,
                .active_state(vasim_50_w_out_9));




/*wire vasim_50_w_out_10;
*/

wire vasim_50_lut_match_10;
wire vasim_50_w_match_10;

    
    
    

LUT_Match_vasim_50_10 #(8) lut_match_vasim_50_10(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_10));


assign vasim_50_w_match_10 = vasim_50_lut_match_10 ;

STE #(.fan_in(1)) vasim_50_ste_10 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_9 }),
                .match(vasim_50_w_match_10) ,
                .active_state(vasim_50_w_out_10));




/*wire vasim_50_w_out_11;
*/

wire vasim_50_lut_match_11;
wire vasim_50_w_match_11;

    
    
    

LUT_Match_vasim_50_11 #(8) lut_match_vasim_50_11(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_11));


assign vasim_50_w_match_11 = vasim_50_lut_match_11 ;

STE #(.fan_in(1)) vasim_50_ste_11 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_10 }),
                .match(vasim_50_w_match_11) ,
                .active_state(vasim_50_w_out_11));




/*wire vasim_50_w_out_12;
*/

wire vasim_50_lut_match_12;
wire vasim_50_w_match_12;

    
    
    

LUT_Match_vasim_50_12 #(8) lut_match_vasim_50_12(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_12));


assign vasim_50_w_match_12 = vasim_50_lut_match_12 ;

STE #(.fan_in(1)) vasim_50_ste_12 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_1 }),
                .match(vasim_50_w_match_12) ,
                .active_state(vasim_50_w_out_12));




/*wire vasim_50_w_out_13;
*/

wire vasim_50_lut_match_13;
wire vasim_50_w_match_13;

    
    
    

LUT_Match_vasim_50_13 #(8) lut_match_vasim_50_13(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_13));


assign vasim_50_w_match_13 = vasim_50_lut_match_13 ;

STE #(.fan_in(1)) vasim_50_ste_13 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_11 }),
                .match(vasim_50_w_match_13) ,
                .active_state(vasim_50_w_out_13));




/*wire vasim_50_w_out_14;
*/

wire vasim_50_lut_match_14;
wire vasim_50_w_match_14;

    
    
    

LUT_Match_vasim_50_14 #(8) lut_match_vasim_50_14(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_14));


assign vasim_50_w_match_14 = vasim_50_lut_match_14 ;

STE #(.fan_in(1)) vasim_50_ste_14 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_13 }),
                .match(vasim_50_w_match_14) ,
                .active_state(vasim_50_w_out_14));




/*wire vasim_50_w_out_15;
*/

wire vasim_50_lut_match_15;
wire vasim_50_w_match_15;

    
    
    

LUT_Match_vasim_50_15 #(8) lut_match_vasim_50_15(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_15));


assign vasim_50_w_match_15 = vasim_50_lut_match_15 ;

STE #(.fan_in(1)) vasim_50_ste_15 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_14 }),
                .match(vasim_50_w_match_15) ,
                .active_state(vasim_50_w_out_15));




/*wire vasim_50_w_out_16;
*/

wire vasim_50_lut_match_16;
wire vasim_50_w_match_16;

    
    
    

LUT_Match_vasim_50_16 #(8) lut_match_vasim_50_16(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_16));


assign vasim_50_w_match_16 = vasim_50_lut_match_16 ;

STE #(.fan_in(1)) vasim_50_ste_16 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_15 }),
                .match(vasim_50_w_match_16) ,
                .active_state(vasim_50_w_out_16));




/*wire vasim_50_w_out_17;
*/

wire vasim_50_lut_match_17;
wire vasim_50_w_match_17;

    
    
    

LUT_Match_vasim_50_17 #(8) lut_match_vasim_50_17(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_17));


assign vasim_50_w_match_17 = vasim_50_lut_match_17 ;

STE #(.fan_in(1)) vasim_50_ste_17 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_16 }),
                .match(vasim_50_w_match_17) ,
                .active_state(vasim_50_w_out_17));




/*wire vasim_50_w_out_18;
*/

wire vasim_50_lut_match_18;
wire vasim_50_w_match_18;

    
    
    

LUT_Match_vasim_50_18 #(8) lut_match_vasim_50_18(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_18));


assign vasim_50_w_match_18 = vasim_50_lut_match_18 ;

STE #(.fan_in(1)) vasim_50_ste_18 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_17 }),
                .match(vasim_50_w_match_18) ,
                .active_state(vasim_50_w_out_18));




/*wire vasim_50_w_out_19;
*/

wire vasim_50_lut_match_19;
wire vasim_50_w_match_19;

    
    
    

LUT_Match_vasim_50_19 #(8) lut_match_vasim_50_19(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_19));


assign vasim_50_w_match_19 = vasim_50_lut_match_19 ;

STE #(.fan_in(1)) vasim_50_ste_19 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_18 }),
                .match(vasim_50_w_match_19) ,
                .active_state(vasim_50_w_out_19));




/*wire vasim_50_w_out_20;
*/

wire vasim_50_lut_match_20;
wire vasim_50_w_match_20;

    
    
    

LUT_Match_vasim_50_20 #(8) lut_match_vasim_50_20(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_20));


assign vasim_50_w_match_20 = vasim_50_lut_match_20 ;

STE #(.fan_in(1)) vasim_50_ste_20 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_19 }),
                .match(vasim_50_w_match_20) ,
                .active_state(vasim_50_w_out_20));




/*wire vasim_50_w_out_21;
*/

wire vasim_50_lut_match_21;
wire vasim_50_w_match_21;

    
    
    

LUT_Match_vasim_50_21 #(8) lut_match_vasim_50_21(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_21));


assign vasim_50_w_match_21 = vasim_50_lut_match_21 ;

STE #(.fan_in(1)) vasim_50_ste_21 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_20 }),
                .match(vasim_50_w_match_21) ,
                .active_state(vasim_50_w_out_21));




/*wire vasim_50_w_out_22;
*/

wire vasim_50_lut_match_22;
wire vasim_50_w_match_22;

    
    
    

LUT_Match_vasim_50_22 #(8) lut_match_vasim_50_22(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_22));


assign vasim_50_w_match_22 = vasim_50_lut_match_22 ;

STE #(.fan_in(1)) vasim_50_ste_22 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_21 }),
                .match(vasim_50_w_match_22) ,
                .active_state(vasim_50_w_out_22));




/*wire vasim_50_w_out_23;
*/

wire vasim_50_lut_match_23;
wire vasim_50_w_match_23;

    
    
    

LUT_Match_vasim_50_23 #(8) lut_match_vasim_50_23(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_23));


assign vasim_50_w_match_23 = vasim_50_lut_match_23 ;

STE #(.fan_in(1)) vasim_50_ste_23 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_12 }),
                .match(vasim_50_w_match_23) ,
                .active_state(vasim_50_w_out_23));




/*wire vasim_50_w_out_24;
*/

wire vasim_50_lut_match_24;
wire vasim_50_w_match_24;

    
    
    

LUT_Match_vasim_50_24 #(8) lut_match_vasim_50_24(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_24));


assign vasim_50_w_match_24 = vasim_50_lut_match_24 ;

STE #(.fan_in(1)) vasim_50_ste_24 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_22 }),
                .match(vasim_50_w_match_24) ,
                .active_state(vasim_50_w_out_24));




/*wire vasim_50_w_out_25;
*/

wire vasim_50_lut_match_25;
wire vasim_50_w_match_25;

    
    
    

LUT_Match_vasim_50_25 #(8) lut_match_vasim_50_25(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_25));


assign vasim_50_w_match_25 = vasim_50_lut_match_25 ;

STE #(.fan_in(1)) vasim_50_ste_25 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_24 }),
                .match(vasim_50_w_match_25) ,
                .active_state(vasim_50_w_out_25));




/*wire vasim_50_w_out_26;
*/

wire vasim_50_lut_match_26;
wire vasim_50_w_match_26;

    
    
    

LUT_Match_vasim_50_26 #(8) lut_match_vasim_50_26(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_26));


assign vasim_50_w_match_26 = vasim_50_lut_match_26 ;

STE #(.fan_in(1)) vasim_50_ste_26 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_25 }),
                .match(vasim_50_w_match_26) ,
                .active_state(vasim_50_w_out_26));




/*wire vasim_50_w_out_27;
*/

wire vasim_50_lut_match_27;
wire vasim_50_w_match_27;

    
    
    

LUT_Match_vasim_50_27 #(8) lut_match_vasim_50_27(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_27));


assign vasim_50_w_match_27 = vasim_50_lut_match_27 ;

STE #(.fan_in(1)) vasim_50_ste_27 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_26 }),
                .match(vasim_50_w_match_27) ,
                .active_state(vasim_50_w_out_27));




/*wire vasim_50_w_out_28;
*/

wire vasim_50_lut_match_28;
wire vasim_50_w_match_28;

    
    
    

LUT_Match_vasim_50_28 #(8) lut_match_vasim_50_28(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_28));


assign vasim_50_w_match_28 = vasim_50_lut_match_28 ;

STE #(.fan_in(1)) vasim_50_ste_28 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_27 }),
                .match(vasim_50_w_match_28) ,
                .active_state(vasim_50_w_out_28));




/*wire vasim_50_w_out_29;
*/

wire vasim_50_lut_match_29;
wire vasim_50_w_match_29;

    
    
    

LUT_Match_vasim_50_29 #(8) lut_match_vasim_50_29(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_29));


assign vasim_50_w_match_29 = vasim_50_lut_match_29 ;

STE #(.fan_in(1)) vasim_50_ste_29 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_28 }),
                .match(vasim_50_w_match_29) ,
                .active_state(vasim_50_w_out_29));




/*wire vasim_50_w_out_30;
*/

wire vasim_50_lut_match_30;
wire vasim_50_w_match_30;

    
    
    

LUT_Match_vasim_50_30 #(8) lut_match_vasim_50_30(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_30));


assign vasim_50_w_match_30 = vasim_50_lut_match_30 ;

STE #(.fan_in(1)) vasim_50_ste_30 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_29 }),
                .match(vasim_50_w_match_30) ,
                .active_state(vasim_50_w_out_30));




/*wire vasim_50_w_out_31;
*/

wire vasim_50_lut_match_31;
wire vasim_50_w_match_31;

    
    
    

LUT_Match_vasim_50_31 #(8) lut_match_vasim_50_31(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_31));


assign vasim_50_w_match_31 = vasim_50_lut_match_31 ;

STE #(.fan_in(1)) vasim_50_ste_31 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_30 }),
                .match(vasim_50_w_match_31) ,
                .active_state(vasim_50_w_out_31));




/*wire vasim_50_w_out_32;
*/

wire vasim_50_lut_match_32;
wire vasim_50_w_match_32;

    
    
    

LUT_Match_vasim_50_32 #(8) lut_match_vasim_50_32(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_32));


assign vasim_50_w_match_32 = vasim_50_lut_match_32 ;

STE #(.fan_in(1)) vasim_50_ste_32 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_31 }),
                .match(vasim_50_w_match_32) ,
                .active_state(vasim_50_w_out_32));




/*wire vasim_50_w_out_33;
*/

wire vasim_50_lut_match_33;
wire vasim_50_w_match_33;

    
    
    

LUT_Match_vasim_50_33 #(8) lut_match_vasim_50_33(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_33));


assign vasim_50_w_match_33 = vasim_50_lut_match_33 ;

STE #(.fan_in(1)) vasim_50_ste_33 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_32 }),
                .match(vasim_50_w_match_33) ,
                .active_state(vasim_50_w_out_33));




/*wire vasim_50_w_out_34;
*/

wire vasim_50_lut_match_34;
wire vasim_50_w_match_34;

    
    
    

LUT_Match_vasim_50_34 #(8) lut_match_vasim_50_34(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_34));


assign vasim_50_w_match_34 = vasim_50_lut_match_34 ;

STE #(.fan_in(1)) vasim_50_ste_34 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_23 }),
                .match(vasim_50_w_match_34) ,
                .active_state(vasim_50_w_out_34));




/*wire vasim_50_w_out_35;
*/

wire vasim_50_lut_match_35;
wire vasim_50_w_match_35;

    
    
    

LUT_Match_vasim_50_35 #(8) lut_match_vasim_50_35(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_35));


assign vasim_50_w_match_35 = vasim_50_lut_match_35 ;

STE #(.fan_in(1)) vasim_50_ste_35 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_33 }),
                .match(vasim_50_w_match_35) ,
                .active_state(vasim_50_w_out_35));




/*wire vasim_50_w_out_36;
*/

wire vasim_50_lut_match_36;
wire vasim_50_w_match_36;

    
    
    

LUT_Match_vasim_50_36 #(8) lut_match_vasim_50_36(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_36));


assign vasim_50_w_match_36 = vasim_50_lut_match_36 ;

STE #(.fan_in(1)) vasim_50_ste_36 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_35 }),
                .match(vasim_50_w_match_36) ,
                .active_state(vasim_50_w_out_36));




/*wire vasim_50_w_out_37;
*/

wire vasim_50_lut_match_37;
wire vasim_50_w_match_37;

    
    
    

LUT_Match_vasim_50_37 #(8) lut_match_vasim_50_37(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_37));


assign vasim_50_w_match_37 = vasim_50_lut_match_37 ;

STE #(.fan_in(1)) vasim_50_ste_37 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_36 }),
                .match(vasim_50_w_match_37) ,
                .active_state(vasim_50_w_out_37));




/*wire vasim_50_w_out_38;
*/

wire vasim_50_lut_match_38;
wire vasim_50_w_match_38;

    
    
    

LUT_Match_vasim_50_38 #(8) lut_match_vasim_50_38(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_38));


assign vasim_50_w_match_38 = vasim_50_lut_match_38 ;

STE #(.fan_in(1)) vasim_50_ste_38 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_37 }),
                .match(vasim_50_w_match_38) ,
                .active_state(vasim_50_w_out_38));




/*wire vasim_50_w_out_39;
*/

wire vasim_50_lut_match_39;
wire vasim_50_w_match_39;

    
    
    

LUT_Match_vasim_50_39 #(8) lut_match_vasim_50_39(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_39));


assign vasim_50_w_match_39 = vasim_50_lut_match_39 ;

STE #(.fan_in(1)) vasim_50_ste_39 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_38 }),
                .match(vasim_50_w_match_39) ,
                .active_state(vasim_50_w_out_39));




/*wire vasim_50_w_out_40;
*/

wire vasim_50_lut_match_40;
wire vasim_50_w_match_40;

    
    
    

LUT_Match_vasim_50_40 #(8) lut_match_vasim_50_40(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_40));


assign vasim_50_w_match_40 = vasim_50_lut_match_40 ;

STE #(.fan_in(1)) vasim_50_ste_40 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_39 }),
                .match(vasim_50_w_match_40) ,
                .active_state(vasim_50_w_out_40));




/*wire vasim_50_w_out_41;
*/

wire vasim_50_lut_match_41;
wire vasim_50_w_match_41;

    
    
    

LUT_Match_vasim_50_41 #(8) lut_match_vasim_50_41(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_41));


assign vasim_50_w_match_41 = vasim_50_lut_match_41 ;

STE #(.fan_in(1)) vasim_50_ste_41 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_40 }),
                .match(vasim_50_w_match_41) ,
                .active_state(vasim_50_w_out_41));




/*wire vasim_50_w_out_42;
*/

wire vasim_50_lut_match_42;
wire vasim_50_w_match_42;

    
    
    

LUT_Match_vasim_50_42 #(8) lut_match_vasim_50_42(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_42));


assign vasim_50_w_match_42 = vasim_50_lut_match_42 ;

STE #(.fan_in(1)) vasim_50_ste_42 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_41 }),
                .match(vasim_50_w_match_42) ,
                .active_state(vasim_50_w_out_42));




/*wire vasim_50_w_out_43;
*/

wire vasim_50_lut_match_43;
wire vasim_50_w_match_43;

    
    
    

LUT_Match_vasim_50_43 #(8) lut_match_vasim_50_43(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_43));


assign vasim_50_w_match_43 = vasim_50_lut_match_43 ;

STE #(.fan_in(1)) vasim_50_ste_43 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_42 }),
                .match(vasim_50_w_match_43) ,
                .active_state(vasim_50_w_out_43));




/*wire vasim_50_w_out_44;
*/

wire vasim_50_lut_match_44;
wire vasim_50_w_match_44;

    
    
    

LUT_Match_vasim_50_44 #(8) lut_match_vasim_50_44(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_44));


assign vasim_50_w_match_44 = vasim_50_lut_match_44 ;

STE #(.fan_in(1)) vasim_50_ste_44 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_43 }),
                .match(vasim_50_w_match_44) ,
                .active_state(vasim_50_w_out_44));




/*wire vasim_50_w_out_45;
*/

wire vasim_50_lut_match_45;
wire vasim_50_w_match_45;

    
    
    

LUT_Match_vasim_50_45 #(8) lut_match_vasim_50_45(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_45));


assign vasim_50_w_match_45 = vasim_50_lut_match_45 ;

STE #(.fan_in(1)) vasim_50_ste_45 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_34 }),
                .match(vasim_50_w_match_45) ,
                .active_state(vasim_50_w_out_45));




/*wire vasim_50_w_out_46;
*/

wire vasim_50_lut_match_46;
wire vasim_50_w_match_46;

    
    
    

LUT_Match_vasim_50_46 #(8) lut_match_vasim_50_46(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_46));


assign vasim_50_w_match_46 = vasim_50_lut_match_46 ;

STE #(.fan_in(1)) vasim_50_ste_46 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_44 }),
                .match(vasim_50_w_match_46) ,
                .active_state(vasim_50_w_out_46));




/*wire vasim_50_w_out_47;
*/

wire vasim_50_lut_match_47;
wire vasim_50_w_match_47;

    
    
    

LUT_Match_vasim_50_47 #(8) lut_match_vasim_50_47(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_47));


assign vasim_50_w_match_47 = vasim_50_lut_match_47 ;

STE #(.fan_in(1)) vasim_50_ste_47 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_46 }),
                .match(vasim_50_w_match_47) ,
                .active_state(vasim_50_w_out_47));




/*wire vasim_50_w_out_48;
*/

wire vasim_50_lut_match_48;
wire vasim_50_w_match_48;

    
    
    

LUT_Match_vasim_50_48 #(8) lut_match_vasim_50_48(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_48));


assign vasim_50_w_match_48 = vasim_50_lut_match_48 ;

STE #(.fan_in(1)) vasim_50_ste_48 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_47 }),
                .match(vasim_50_w_match_48) ,
                .active_state(vasim_50_w_out_48));




/*wire vasim_50_w_out_49;
*/

wire vasim_50_lut_match_49;
wire vasim_50_w_match_49;

    
    
    

LUT_Match_vasim_50_49 #(8) lut_match_vasim_50_49(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_49));


assign vasim_50_w_match_49 = vasim_50_lut_match_49 ;

STE #(.fan_in(1)) vasim_50_ste_49 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_48 }),
                .match(vasim_50_w_match_49) ,
                .active_state(vasim_50_w_out_49));




/*wire vasim_50_w_out_50;
*/

wire vasim_50_lut_match_50;
wire vasim_50_w_match_50;

    
    
    

LUT_Match_vasim_50_50 #(8) lut_match_vasim_50_50(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_50));


assign vasim_50_w_match_50 = vasim_50_lut_match_50 ;

STE #(.fan_in(1)) vasim_50_ste_50 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_49 }),
                .match(vasim_50_w_match_50) ,
                .active_state(vasim_50_w_out_50));




/*wire vasim_50_w_out_51;
*/

wire vasim_50_lut_match_51;
wire vasim_50_w_match_51;

    
    
    

LUT_Match_vasim_50_51 #(8) lut_match_vasim_50_51(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_51));


assign vasim_50_w_match_51 = vasim_50_lut_match_51 ;

STE #(.fan_in(1)) vasim_50_ste_51 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_50 }),
                .match(vasim_50_w_match_51) ,
                .active_state(vasim_50_w_out_51));




/*wire vasim_50_w_out_52;
*/

wire vasim_50_lut_match_52;
wire vasim_50_w_match_52;

    
    
    

LUT_Match_vasim_50_52 #(8) lut_match_vasim_50_52(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_52));


assign vasim_50_w_match_52 = vasim_50_lut_match_52 ;

STE #(.fan_in(1)) vasim_50_ste_52 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_51 }),
                .match(vasim_50_w_match_52) ,
                .active_state(vasim_50_w_out_52));




/*wire vasim_50_w_out_53;
*/

wire vasim_50_lut_match_53;
wire vasim_50_w_match_53;

    
    
    

LUT_Match_vasim_50_53 #(8) lut_match_vasim_50_53(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_53));


assign vasim_50_w_match_53 = vasim_50_lut_match_53 ;

STE #(.fan_in(1)) vasim_50_ste_53 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_52 }),
                .match(vasim_50_w_match_53) ,
                .active_state(vasim_50_w_out_53));




/*wire vasim_50_w_out_54;
*/

wire vasim_50_lut_match_54;
wire vasim_50_w_match_54;

    
    
    

LUT_Match_vasim_50_54 #(8) lut_match_vasim_50_54(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_54));


assign vasim_50_w_match_54 = vasim_50_lut_match_54 ;

STE #(.fan_in(1)) vasim_50_ste_54 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_53 }),
                .match(vasim_50_w_match_54) ,
                .active_state(vasim_50_w_out_54));




/*wire vasim_50_w_out_55;
*/

wire vasim_50_lut_match_55;
wire vasim_50_w_match_55;

    
    
    

LUT_Match_vasim_50_55 #(8) lut_match_vasim_50_55(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_55));


assign vasim_50_w_match_55 = vasim_50_lut_match_55 ;

STE #(.fan_in(1)) vasim_50_ste_55 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_54 }),
                .match(vasim_50_w_match_55) ,
                .active_state(vasim_50_w_out_55));




/*wire vasim_50_w_out_56;
*/

wire vasim_50_lut_match_56;
wire vasim_50_w_match_56;

    
    
    

LUT_Match_vasim_50_56 #(8) lut_match_vasim_50_56(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_56));


assign vasim_50_w_match_56 = vasim_50_lut_match_56 ;

STE #(.fan_in(1)) vasim_50_ste_56 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_45 }),
                .match(vasim_50_w_match_56) ,
                .active_state(vasim_50_w_out_56));




/*wire vasim_50_w_out_57;
*/

wire vasim_50_lut_match_57;
wire vasim_50_w_match_57;

    
    
    

LUT_Match_vasim_50_57 #(8) lut_match_vasim_50_57(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_57));


assign vasim_50_w_match_57 = vasim_50_lut_match_57 ;

STE #(.fan_in(1)) vasim_50_ste_57 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_55 }),
                .match(vasim_50_w_match_57) ,
                .active_state(vasim_50_w_out_57));




/*wire vasim_50_w_out_58;
*/

wire vasim_50_lut_match_58;
wire vasim_50_w_match_58;

    
    
    

LUT_Match_vasim_50_58 #(8) lut_match_vasim_50_58(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_58));


assign vasim_50_w_match_58 = vasim_50_lut_match_58 ;

STE #(.fan_in(1)) vasim_50_ste_58 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_57 }),
                .match(vasim_50_w_match_58) ,
                .active_state(vasim_50_w_out_58));




/*wire vasim_50_w_out_59;
*/

wire vasim_50_lut_match_59;
wire vasim_50_w_match_59;

    
    
    

LUT_Match_vasim_50_59 #(8) lut_match_vasim_50_59(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_59));


assign vasim_50_w_match_59 = vasim_50_lut_match_59 ;

STE #(.fan_in(1)) vasim_50_ste_59 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_58 }),
                .match(vasim_50_w_match_59) ,
                .active_state(vasim_50_w_out_59));




/*wire vasim_50_w_out_60;
*/

wire vasim_50_lut_match_60;
wire vasim_50_w_match_60;

    
    
    

LUT_Match_vasim_50_60 #(8) lut_match_vasim_50_60(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_60));


assign vasim_50_w_match_60 = vasim_50_lut_match_60 ;

STE #(.fan_in(1)) vasim_50_ste_60 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_59 }),
                .match(vasim_50_w_match_60) ,
                .active_state(vasim_50_w_out_60));




/*wire vasim_50_w_out_61;
*/

wire vasim_50_lut_match_61;
wire vasim_50_w_match_61;

    
    
    

LUT_Match_vasim_50_61 #(8) lut_match_vasim_50_61(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_61));


assign vasim_50_w_match_61 = vasim_50_lut_match_61 ;

STE #(.fan_in(1)) vasim_50_ste_61 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_60 }),
                .match(vasim_50_w_match_61) ,
                .active_state(vasim_50_w_out_61));




/*wire vasim_50_w_out_62;
*/

wire vasim_50_lut_match_62;
wire vasim_50_w_match_62;

    
    
    

LUT_Match_vasim_50_62 #(8) lut_match_vasim_50_62(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_62));


assign vasim_50_w_match_62 = vasim_50_lut_match_62 ;

STE #(.fan_in(1)) vasim_50_ste_62 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_61 }),
                .match(vasim_50_w_match_62) ,
                .active_state(vasim_50_w_out_62));




/*wire vasim_50_w_out_63;
*/

wire vasim_50_lut_match_63;
wire vasim_50_w_match_63;

    
    
    

LUT_Match_vasim_50_63 #(8) lut_match_vasim_50_63(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_63));


assign vasim_50_w_match_63 = vasim_50_lut_match_63 ;

STE #(.fan_in(1)) vasim_50_ste_63 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_62 }),
                .match(vasim_50_w_match_63) ,
                .active_state(vasim_50_w_out_63));




/*wire vasim_50_w_out_64;
*/

wire vasim_50_lut_match_64;
wire vasim_50_w_match_64;

    
    
    

LUT_Match_vasim_50_64 #(8) lut_match_vasim_50_64(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_64));


assign vasim_50_w_match_64 = vasim_50_lut_match_64 ;

STE #(.fan_in(1)) vasim_50_ste_64 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_63 }),
                .match(vasim_50_w_match_64) ,
                .active_state(vasim_50_w_out_64));




/*wire vasim_50_w_out_65;
*/

wire vasim_50_lut_match_65;
wire vasim_50_w_match_65;

    
    
    

LUT_Match_vasim_50_65 #(8) lut_match_vasim_50_65(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_65));


assign vasim_50_w_match_65 = vasim_50_lut_match_65 ;

STE #(.fan_in(1)) vasim_50_ste_65 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_64 }),
                .match(vasim_50_w_match_65) ,
                .active_state(vasim_50_w_out_65));




/*wire vasim_50_w_out_66;
*/

wire vasim_50_lut_match_66;
wire vasim_50_w_match_66;

    
    
    

LUT_Match_vasim_50_66 #(8) lut_match_vasim_50_66(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_66));


assign vasim_50_w_match_66 = vasim_50_lut_match_66 ;

STE #(.fan_in(1)) vasim_50_ste_66 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_65 }),
                .match(vasim_50_w_match_66) ,
                .active_state(vasim_50_w_out_66));




/*wire vasim_50_w_out_67;
*/

wire vasim_50_lut_match_67;
wire vasim_50_w_match_67;

    
    
    

LUT_Match_vasim_50_67 #(8) lut_match_vasim_50_67(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_67));


assign vasim_50_w_match_67 = vasim_50_lut_match_67 ;

STE #(.fan_in(1)) vasim_50_ste_67 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_56 }),
                .match(vasim_50_w_match_67) ,
                .active_state(vasim_50_w_out_67));




/*wire vasim_50_w_out_68;
*/

wire vasim_50_lut_match_68;
wire vasim_50_w_match_68;

    
    
    

LUT_Match_vasim_50_68 #(8) lut_match_vasim_50_68(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_68));


assign vasim_50_w_match_68 = vasim_50_lut_match_68 ;

STE #(.fan_in(1)) vasim_50_ste_68 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_66 }),
                .match(vasim_50_w_match_68) ,
                .active_state(vasim_50_w_out_68));




/*wire vasim_50_w_out_69;
*/

wire vasim_50_lut_match_69;
wire vasim_50_w_match_69;

    
    
    

LUT_Match_vasim_50_69 #(8) lut_match_vasim_50_69(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_69));


assign vasim_50_w_match_69 = vasim_50_lut_match_69 ;

STE #(.fan_in(1)) vasim_50_ste_69 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_68 }),
                .match(vasim_50_w_match_69) ,
                .active_state(vasim_50_w_out_69));




/*wire vasim_50_w_out_70;
*/

wire vasim_50_lut_match_70;
wire vasim_50_w_match_70;

    
    
    

LUT_Match_vasim_50_70 #(8) lut_match_vasim_50_70(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_70));


assign vasim_50_w_match_70 = vasim_50_lut_match_70 ;

STE #(.fan_in(1)) vasim_50_ste_70 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_69 }),
                .match(vasim_50_w_match_70) ,
                .active_state(vasim_50_w_out_70));




/*wire vasim_50_w_out_71;
*/

wire vasim_50_lut_match_71;
wire vasim_50_w_match_71;

    
    
    

LUT_Match_vasim_50_71 #(8) lut_match_vasim_50_71(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_71));


assign vasim_50_w_match_71 = vasim_50_lut_match_71 ;

STE #(.fan_in(1)) vasim_50_ste_71 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_70 }),
                .match(vasim_50_w_match_71) ,
                .active_state(vasim_50_w_out_71));




/*wire vasim_50_w_out_72;
*/

wire vasim_50_lut_match_72;
wire vasim_50_w_match_72;

    
    
    

LUT_Match_vasim_50_72 #(8) lut_match_vasim_50_72(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_72));


assign vasim_50_w_match_72 = vasim_50_lut_match_72 ;

STE #(.fan_in(1)) vasim_50_ste_72 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_71 }),
                .match(vasim_50_w_match_72) ,
                .active_state(vasim_50_w_out_72));




/*wire vasim_50_w_out_73;
*/

wire vasim_50_lut_match_73;
wire vasim_50_w_match_73;

    
    
    

LUT_Match_vasim_50_73 #(8) lut_match_vasim_50_73(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_73));


assign vasim_50_w_match_73 = vasim_50_lut_match_73 ;

STE #(.fan_in(1)) vasim_50_ste_73 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_72 }),
                .match(vasim_50_w_match_73) ,
                .active_state(vasim_50_w_out_73));




/*wire vasim_50_w_out_74;
*/

wire vasim_50_lut_match_74;
wire vasim_50_w_match_74;

    
    
    

LUT_Match_vasim_50_74 #(8) lut_match_vasim_50_74(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_74));


assign vasim_50_w_match_74 = vasim_50_lut_match_74 ;

STE #(.fan_in(1)) vasim_50_ste_74 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_73 }),
                .match(vasim_50_w_match_74) ,
                .active_state(vasim_50_w_out_74));




/*wire vasim_50_w_out_75;
*/

wire vasim_50_lut_match_75;
wire vasim_50_w_match_75;

    
    
    

LUT_Match_vasim_50_75 #(8) lut_match_vasim_50_75(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_75));


assign vasim_50_w_match_75 = vasim_50_lut_match_75 ;

STE #(.fan_in(1)) vasim_50_ste_75 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_74 }),
                .match(vasim_50_w_match_75) ,
                .active_state(vasim_50_w_out_75));




/*wire vasim_50_w_out_76;
*/

wire vasim_50_lut_match_76;
wire vasim_50_w_match_76;

    
    
    

LUT_Match_vasim_50_76 #(8) lut_match_vasim_50_76(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_76));


assign vasim_50_w_match_76 = vasim_50_lut_match_76 ;

STE #(.fan_in(1)) vasim_50_ste_76 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_75 }),
                .match(vasim_50_w_match_76) ,
                .active_state(vasim_50_w_out_76));




/*wire vasim_50_w_out_77;
*/

wire vasim_50_lut_match_77;
wire vasim_50_w_match_77;

    
    
    

LUT_Match_vasim_50_77 #(8) lut_match_vasim_50_77(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_77));


assign vasim_50_w_match_77 = vasim_50_lut_match_77 ;

STE #(.fan_in(1)) vasim_50_ste_77 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_76 }),
                .match(vasim_50_w_match_77) ,
                .active_state(vasim_50_w_out_77));




/*wire vasim_50_w_out_78;
*/

wire vasim_50_lut_match_78;
wire vasim_50_w_match_78;

    
    
    

LUT_Match_vasim_50_78 #(8) lut_match_vasim_50_78(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_78));


assign vasim_50_w_match_78 = vasim_50_lut_match_78 ;

STE #(.fan_in(1)) vasim_50_ste_78 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_67 }),
                .match(vasim_50_w_match_78) ,
                .active_state(vasim_50_w_out_78));




/*wire vasim_50_w_out_79;
*/

wire vasim_50_lut_match_79;
wire vasim_50_w_match_79;

    
    
    

LUT_Match_vasim_50_79 #(8) lut_match_vasim_50_79(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_79));


assign vasim_50_w_match_79 = vasim_50_lut_match_79 ;

STE #(.fan_in(1)) vasim_50_ste_79 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_77 }),
                .match(vasim_50_w_match_79) ,
                .active_state(vasim_50_w_out_79));




/*wire vasim_50_w_out_80;
*/

wire vasim_50_lut_match_80;
wire vasim_50_w_match_80;

    
    
    

LUT_Match_vasim_50_80 #(8) lut_match_vasim_50_80(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_80));


assign vasim_50_w_match_80 = vasim_50_lut_match_80 ;

STE #(.fan_in(1)) vasim_50_ste_80 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_79 }),
                .match(vasim_50_w_match_80) ,
                .active_state(vasim_50_w_out_80));




/*wire vasim_50_w_out_81;
*/

wire vasim_50_lut_match_81;
wire vasim_50_w_match_81;

    
    
    

LUT_Match_vasim_50_81 #(8) lut_match_vasim_50_81(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_81));


assign vasim_50_w_match_81 = vasim_50_lut_match_81 ;

STE #(.fan_in(1)) vasim_50_ste_81 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_80 }),
                .match(vasim_50_w_match_81) ,
                .active_state(vasim_50_w_out_81));




/*wire vasim_50_w_out_82;
*/

wire vasim_50_lut_match_82;
wire vasim_50_w_match_82;

    
    
    

LUT_Match_vasim_50_82 #(8) lut_match_vasim_50_82(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_82));


assign vasim_50_w_match_82 = vasim_50_lut_match_82 ;

STE #(.fan_in(1)) vasim_50_ste_82 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_81 }),
                .match(vasim_50_w_match_82) ,
                .active_state(vasim_50_w_out_82));




/*wire vasim_50_w_out_83;
*/

wire vasim_50_lut_match_83;
wire vasim_50_w_match_83;

    
    
    

LUT_Match_vasim_50_83 #(8) lut_match_vasim_50_83(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_83));


assign vasim_50_w_match_83 = vasim_50_lut_match_83 ;

STE #(.fan_in(1)) vasim_50_ste_83 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_82 }),
                .match(vasim_50_w_match_83) ,
                .active_state(vasim_50_w_out_83));




/*wire vasim_50_w_out_84;
*/

wire vasim_50_lut_match_84;
wire vasim_50_w_match_84;

    
    
    

LUT_Match_vasim_50_84 #(8) lut_match_vasim_50_84(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_84));


assign vasim_50_w_match_84 = vasim_50_lut_match_84 ;

STE #(.fan_in(1)) vasim_50_ste_84 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_83 }),
                .match(vasim_50_w_match_84) ,
                .active_state(vasim_50_w_out_84));




/*wire vasim_50_w_out_85;
*/

wire vasim_50_lut_match_85;
wire vasim_50_w_match_85;

    
    
    

LUT_Match_vasim_50_85 #(8) lut_match_vasim_50_85(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_85));


assign vasim_50_w_match_85 = vasim_50_lut_match_85 ;

STE #(.fan_in(1)) vasim_50_ste_85 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_84 }),
                .match(vasim_50_w_match_85) ,
                .active_state(vasim_50_w_out_85));




/*wire vasim_50_w_out_86;
*/

wire vasim_50_lut_match_86;
wire vasim_50_w_match_86;

    
    
    

LUT_Match_vasim_50_86 #(8) lut_match_vasim_50_86(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_86));


assign vasim_50_w_match_86 = vasim_50_lut_match_86 ;

STE #(.fan_in(1)) vasim_50_ste_86 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_85 }),
                .match(vasim_50_w_match_86) ,
                .active_state(vasim_50_w_out_86));




/*wire vasim_50_w_out_87;
*/

wire vasim_50_lut_match_87;
wire vasim_50_w_match_87;

    
    
    

LUT_Match_vasim_50_87 #(8) lut_match_vasim_50_87(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_87));


assign vasim_50_w_match_87 = vasim_50_lut_match_87 ;

STE #(.fan_in(1)) vasim_50_ste_87 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_86 }),
                .match(vasim_50_w_match_87) ,
                .active_state(vasim_50_w_out_87));




/*wire vasim_50_w_out_88;
*/

wire vasim_50_lut_match_88;
wire vasim_50_w_match_88;

    
    
    

LUT_Match_vasim_50_88 #(8) lut_match_vasim_50_88(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_88));


assign vasim_50_w_match_88 = vasim_50_lut_match_88 ;

STE #(.fan_in(1)) vasim_50_ste_88 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_87 }),
                .match(vasim_50_w_match_88) ,
                .active_state(vasim_50_w_out_88));




/*wire vasim_50_w_out_89;
*/

wire vasim_50_lut_match_89;
wire vasim_50_w_match_89;

    
    
    

LUT_Match_vasim_50_89 #(8) lut_match_vasim_50_89(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_89));


assign vasim_50_w_match_89 = vasim_50_lut_match_89 ;

STE #(.fan_in(1)) vasim_50_ste_89 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_78 }),
                .match(vasim_50_w_match_89) ,
                .active_state(vasim_50_w_out_89));




/*wire vasim_50_w_out_90;
*/

wire vasim_50_lut_match_90;
wire vasim_50_w_match_90;

    
    
    

LUT_Match_vasim_50_90 #(8) lut_match_vasim_50_90(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_90));


assign vasim_50_w_match_90 = vasim_50_lut_match_90 ;

STE #(.fan_in(1)) vasim_50_ste_90 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_88 }),
                .match(vasim_50_w_match_90) ,
                .active_state(vasim_50_w_out_90));




/*wire vasim_50_w_out_91;
*/

wire vasim_50_lut_match_91;
wire vasim_50_w_match_91;

    
    
    

LUT_Match_vasim_50_91 #(8) lut_match_vasim_50_91(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_91));


assign vasim_50_w_match_91 = vasim_50_lut_match_91 ;

STE #(.fan_in(1)) vasim_50_ste_91 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_90 }),
                .match(vasim_50_w_match_91) ,
                .active_state(vasim_50_w_out_91));




/*wire vasim_50_w_out_92;
*/

wire vasim_50_lut_match_92;
wire vasim_50_w_match_92;

    
    
    

LUT_Match_vasim_50_92 #(8) lut_match_vasim_50_92(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_92));


assign vasim_50_w_match_92 = vasim_50_lut_match_92 ;

STE #(.fan_in(1)) vasim_50_ste_92 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_91 }),
                .match(vasim_50_w_match_92) ,
                .active_state(vasim_50_w_out_92));




/*wire vasim_50_w_out_93;
*/

wire vasim_50_lut_match_93;
wire vasim_50_w_match_93;

    
    
    

LUT_Match_vasim_50_93 #(8) lut_match_vasim_50_93(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_93));


assign vasim_50_w_match_93 = vasim_50_lut_match_93 ;

STE #(.fan_in(1)) vasim_50_ste_93 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_92 }),
                .match(vasim_50_w_match_93) ,
                .active_state(vasim_50_w_out_93));




/*wire vasim_50_w_out_94;
*/

wire vasim_50_lut_match_94;
wire vasim_50_w_match_94;

    
    
    

LUT_Match_vasim_50_94 #(8) lut_match_vasim_50_94(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_94));


assign vasim_50_w_match_94 = vasim_50_lut_match_94 ;

STE #(.fan_in(1)) vasim_50_ste_94 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_93 }),
                .match(vasim_50_w_match_94) ,
                .active_state(vasim_50_w_out_94));




/*wire vasim_50_w_out_95;
*/

wire vasim_50_lut_match_95;
wire vasim_50_w_match_95;

    
    
    

LUT_Match_vasim_50_95 #(8) lut_match_vasim_50_95(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_95));


assign vasim_50_w_match_95 = vasim_50_lut_match_95 ;

STE #(.fan_in(1)) vasim_50_ste_95 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_94 }),
                .match(vasim_50_w_match_95) ,
                .active_state(vasim_50_w_out_95));




/*wire vasim_50_w_out_96;
*/

wire vasim_50_lut_match_96;
wire vasim_50_w_match_96;

    
    
    

LUT_Match_vasim_50_96 #(8) lut_match_vasim_50_96(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_96));


assign vasim_50_w_match_96 = vasim_50_lut_match_96 ;

STE #(.fan_in(1)) vasim_50_ste_96 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_95 }),
                .match(vasim_50_w_match_96) ,
                .active_state(vasim_50_w_out_96));




/*wire vasim_50_w_out_97;
*/

wire vasim_50_lut_match_97;
wire vasim_50_w_match_97;

    
    
    

LUT_Match_vasim_50_97 #(8) lut_match_vasim_50_97(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_97));


assign vasim_50_w_match_97 = vasim_50_lut_match_97 ;

STE #(.fan_in(1)) vasim_50_ste_97 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_96 }),
                .match(vasim_50_w_match_97) ,
                .active_state(vasim_50_w_out_97));




/*wire vasim_50_w_out_98;
*/

wire vasim_50_lut_match_98;
wire vasim_50_w_match_98;

    
    
    

LUT_Match_vasim_50_98 #(8) lut_match_vasim_50_98(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_98));


assign vasim_50_w_match_98 = vasim_50_lut_match_98 ;

STE #(.fan_in(1)) vasim_50_ste_98 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_97 }),
                .match(vasim_50_w_match_98) ,
                .active_state(vasim_50_w_out_98));




/*wire vasim_50_w_out_99;
*/

wire vasim_50_lut_match_99;
wire vasim_50_w_match_99;

    
    
    

LUT_Match_vasim_50_99 #(8) lut_match_vasim_50_99(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_99));


assign vasim_50_w_match_99 = vasim_50_lut_match_99 ;

STE #(.fan_in(1)) vasim_50_ste_99 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_98 }),
                .match(vasim_50_w_match_99) ,
                .active_state(vasim_50_w_out_99));




/*wire vasim_50_w_out_100;
*/

wire vasim_50_lut_match_100;
wire vasim_50_w_match_100;

    
    
    

LUT_Match_vasim_50_100 #(8) lut_match_vasim_50_100(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_100));


assign vasim_50_w_match_100 = vasim_50_lut_match_100 ;

STE #(.fan_in(1)) vasim_50_ste_100 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_89 }),
                .match(vasim_50_w_match_100) ,
                .active_state(vasim_50_w_out_100));




/*wire vasim_50_w_out_101;
*/

wire vasim_50_lut_match_101;
wire vasim_50_w_match_101;

    
    
    

LUT_Match_vasim_50_101 #(8) lut_match_vasim_50_101(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_101));


assign vasim_50_w_match_101 = vasim_50_lut_match_101 ;

STE #(.fan_in(1)) vasim_50_ste_101 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_99 }),
                .match(vasim_50_w_match_101) ,
                .active_state(vasim_50_w_out_101));




/*wire vasim_50_w_out_102;
*/

wire vasim_50_lut_match_102;
wire vasim_50_w_match_102;

    
    
    

LUT_Match_vasim_50_102 #(8) lut_match_vasim_50_102(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_102));


assign vasim_50_w_match_102 = vasim_50_lut_match_102 ;

STE #(.fan_in(1)) vasim_50_ste_102 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_101 }),
                .match(vasim_50_w_match_102) ,
                .active_state(vasim_50_w_out_102));




/*wire vasim_50_w_out_103;
*/

wire vasim_50_lut_match_103;
wire vasim_50_w_match_103;

    
    
    

LUT_Match_vasim_50_103 #(8) lut_match_vasim_50_103(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_103));


assign vasim_50_w_match_103 = vasim_50_lut_match_103 ;

STE #(.fan_in(1)) vasim_50_ste_103 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_102 }),
                .match(vasim_50_w_match_103) ,
                .active_state(vasim_50_w_out_103));




/*wire vasim_50_w_out_104;
*/

wire vasim_50_lut_match_104;
wire vasim_50_w_match_104;

    
    
    

LUT_Match_vasim_50_104 #(8) lut_match_vasim_50_104(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_104));


assign vasim_50_w_match_104 = vasim_50_lut_match_104 ;

STE #(.fan_in(1)) vasim_50_ste_104 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_103 }),
                .match(vasim_50_w_match_104) ,
                .active_state(vasim_50_w_out_104));




/*wire vasim_50_w_out_105;
*/

wire vasim_50_lut_match_105;
wire vasim_50_w_match_105;

    
    
    

LUT_Match_vasim_50_105 #(8) lut_match_vasim_50_105(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_105));


assign vasim_50_w_match_105 = vasim_50_lut_match_105 ;

STE #(.fan_in(1)) vasim_50_ste_105 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_104 }),
                .match(vasim_50_w_match_105) ,
                .active_state(vasim_50_w_out_105));




/*wire vasim_50_w_out_106;
*/

wire vasim_50_lut_match_106;
wire vasim_50_w_match_106;

    
    
    

LUT_Match_vasim_50_106 #(8) lut_match_vasim_50_106(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_106));


assign vasim_50_w_match_106 = vasim_50_lut_match_106 ;

STE #(.fan_in(1)) vasim_50_ste_106 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_105 }),
                .match(vasim_50_w_match_106) ,
                .active_state(vasim_50_w_out_106));




/*wire vasim_50_w_out_107;
*/

wire vasim_50_lut_match_107;
wire vasim_50_w_match_107;

    
    
    

LUT_Match_vasim_50_107 #(8) lut_match_vasim_50_107(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_107));


assign vasim_50_w_match_107 = vasim_50_lut_match_107 ;

STE #(.fan_in(1)) vasim_50_ste_107 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_106 }),
                .match(vasim_50_w_match_107) ,
                .active_state(vasim_50_w_out_107));




/*wire vasim_50_w_out_108;
*/

wire vasim_50_lut_match_108;
wire vasim_50_w_match_108;

    
    
    

LUT_Match_vasim_50_108 #(8) lut_match_vasim_50_108(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_108));


assign vasim_50_w_match_108 = vasim_50_lut_match_108 ;

STE #(.fan_in(1)) vasim_50_ste_108 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_107 }),
                .match(vasim_50_w_match_108) ,
                .active_state(vasim_50_w_out_108));




/*wire vasim_50_w_out_109;
*/

wire vasim_50_lut_match_109;
wire vasim_50_w_match_109;

    
    
    

LUT_Match_vasim_50_109 #(8) lut_match_vasim_50_109(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_109));


assign vasim_50_w_match_109 = vasim_50_lut_match_109 ;

STE #(.fan_in(1)) vasim_50_ste_109 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_108 }),
                .match(vasim_50_w_match_109) ,
                .active_state(vasim_50_w_out_109));




/*wire vasim_50_w_out_110;
*/

wire vasim_50_lut_match_110;
wire vasim_50_w_match_110;

    
    
    

LUT_Match_vasim_50_110 #(8) lut_match_vasim_50_110(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_110));


assign vasim_50_w_match_110 = vasim_50_lut_match_110 ;

STE #(.fan_in(1)) vasim_50_ste_110 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_109 }),
                .match(vasim_50_w_match_110) ,
                .active_state(vasim_50_w_out_110));




/*wire vasim_50_w_out_111;
*/

wire vasim_50_lut_match_111;
wire vasim_50_w_match_111;

    
    
    

LUT_Match_vasim_50_111 #(8) lut_match_vasim_50_111(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_111));


assign vasim_50_w_match_111 = vasim_50_lut_match_111 ;

STE #(.fan_in(1)) vasim_50_ste_111 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_100 }),
                .match(vasim_50_w_match_111) ,
                .active_state(vasim_50_w_out_111));




/*wire vasim_50_w_out_112;
*/

wire vasim_50_lut_match_112;
wire vasim_50_w_match_112;

    
    
    

LUT_Match_vasim_50_112 #(8) lut_match_vasim_50_112(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_112));


assign vasim_50_w_match_112 = vasim_50_lut_match_112 ;

STE #(.fan_in(1)) vasim_50_ste_112 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_110 }),
                .match(vasim_50_w_match_112) ,
                .active_state(vasim_50_w_out_112));




/*wire vasim_50_w_out_113;
*/

wire vasim_50_lut_match_113;
wire vasim_50_w_match_113;

    
    
    

LUT_Match_vasim_50_113 #(8) lut_match_vasim_50_113(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_113));


assign vasim_50_w_match_113 = vasim_50_lut_match_113 ;

STE #(.fan_in(1)) vasim_50_ste_113 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_112 }),
                .match(vasim_50_w_match_113) ,
                .active_state(vasim_50_w_out_113));




/*wire vasim_50_w_out_114;
*/

wire vasim_50_lut_match_114;
wire vasim_50_w_match_114;

    
    
    

LUT_Match_vasim_50_114 #(8) lut_match_vasim_50_114(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_114));


assign vasim_50_w_match_114 = vasim_50_lut_match_114 ;

STE #(.fan_in(1)) vasim_50_ste_114 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_113 }),
                .match(vasim_50_w_match_114) ,
                .active_state(vasim_50_w_out_114));




/*wire vasim_50_w_out_115;
*/

wire vasim_50_lut_match_115;
wire vasim_50_w_match_115;

    
    
    

LUT_Match_vasim_50_115 #(8) lut_match_vasim_50_115(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_115));


assign vasim_50_w_match_115 = vasim_50_lut_match_115 ;

STE #(.fan_in(1)) vasim_50_ste_115 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_114 }),
                .match(vasim_50_w_match_115) ,
                .active_state(vasim_50_w_out_115));




/*wire vasim_50_w_out_116;
*/

wire vasim_50_lut_match_116;
wire vasim_50_w_match_116;

    
    
    

LUT_Match_vasim_50_116 #(8) lut_match_vasim_50_116(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_116));


assign vasim_50_w_match_116 = vasim_50_lut_match_116 ;

STE #(.fan_in(1)) vasim_50_ste_116 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_115 }),
                .match(vasim_50_w_match_116) ,
                .active_state(vasim_50_w_out_116));




/*wire vasim_50_w_out_117;
*/

wire vasim_50_lut_match_117;
wire vasim_50_w_match_117;

    
    
    

LUT_Match_vasim_50_117 #(8) lut_match_vasim_50_117(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_117));


assign vasim_50_w_match_117 = vasim_50_lut_match_117 ;

STE #(.fan_in(1)) vasim_50_ste_117 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_116 }),
                .match(vasim_50_w_match_117) ,
                .active_state(vasim_50_w_out_117));




/*wire vasim_50_w_out_118;
*/

wire vasim_50_lut_match_118;
wire vasim_50_w_match_118;

    
    
    

LUT_Match_vasim_50_118 #(8) lut_match_vasim_50_118(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_118));


assign vasim_50_w_match_118 = vasim_50_lut_match_118 ;

STE #(.fan_in(1)) vasim_50_ste_118 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_117 }),
                .match(vasim_50_w_match_118) ,
                .active_state(vasim_50_w_out_118));




/*wire vasim_50_w_out_119;
*/

wire vasim_50_lut_match_119;
wire vasim_50_w_match_119;

    
    
    

LUT_Match_vasim_50_119 #(8) lut_match_vasim_50_119(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_119));


assign vasim_50_w_match_119 = vasim_50_lut_match_119 ;

STE #(.fan_in(1)) vasim_50_ste_119 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_118 }),
                .match(vasim_50_w_match_119) ,
                .active_state(vasim_50_w_out_119));




/*wire vasim_50_w_out_120;
*/

wire vasim_50_lut_match_120;
wire vasim_50_w_match_120;

    
    
    

LUT_Match_vasim_50_120 #(8) lut_match_vasim_50_120(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_120));


assign vasim_50_w_match_120 = vasim_50_lut_match_120 ;

STE #(.fan_in(1)) vasim_50_ste_120 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_119 }),
                .match(vasim_50_w_match_120) ,
                .active_state(vasim_50_w_out_120));




/*wire vasim_50_w_out_121;
*/

wire vasim_50_lut_match_121;
wire vasim_50_w_match_121;

    
    
    

LUT_Match_vasim_50_121 #(8) lut_match_vasim_50_121(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_121));


assign vasim_50_w_match_121 = vasim_50_lut_match_121 ;

STE #(.fan_in(1)) vasim_50_ste_121 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_120 }),
                .match(vasim_50_w_match_121) ,
                .active_state(vasim_50_w_out_121));




/*wire vasim_50_w_out_122;
*/

wire vasim_50_lut_match_122;
wire vasim_50_w_match_122;

    
    
    

LUT_Match_vasim_50_122 #(8) lut_match_vasim_50_122(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_122));


assign vasim_50_w_match_122 = vasim_50_lut_match_122 ;

STE #(.fan_in(1)) vasim_50_ste_122 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_111 }),
                .match(vasim_50_w_match_122) ,
                .active_state(vasim_50_w_out_122));




/*wire vasim_50_w_out_123;
*/

wire vasim_50_lut_match_123;
wire vasim_50_w_match_123;

    
    
    

LUT_Match_vasim_50_123 #(8) lut_match_vasim_50_123(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_123));


assign vasim_50_w_match_123 = vasim_50_lut_match_123 ;

STE #(.fan_in(1)) vasim_50_ste_123 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_121 }),
                .match(vasim_50_w_match_123) ,
                .active_state(vasim_50_w_out_123));




/*wire vasim_50_w_out_124;
*/

wire vasim_50_lut_match_124;
wire vasim_50_w_match_124;

    
    
    

LUT_Match_vasim_50_124 #(8) lut_match_vasim_50_124(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_124));


assign vasim_50_w_match_124 = vasim_50_lut_match_124 ;

STE #(.fan_in(1)) vasim_50_ste_124 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_123 }),
                .match(vasim_50_w_match_124) ,
                .active_state(vasim_50_w_out_124));




/*wire vasim_50_w_out_125;
*/

wire vasim_50_lut_match_125;
wire vasim_50_w_match_125;

    
    
    

LUT_Match_vasim_50_125 #(8) lut_match_vasim_50_125(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_125));


assign vasim_50_w_match_125 = vasim_50_lut_match_125 ;

STE #(.fan_in(1)) vasim_50_ste_125 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_124 }),
                .match(vasim_50_w_match_125) ,
                .active_state(vasim_50_w_out_125));




/*wire vasim_50_w_out_126;
*/

wire vasim_50_lut_match_126;
wire vasim_50_w_match_126;

    
    
    

LUT_Match_vasim_50_126 #(8) lut_match_vasim_50_126(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_126));


assign vasim_50_w_match_126 = vasim_50_lut_match_126 ;

STE #(.fan_in(1)) vasim_50_ste_126 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_125 }),
                .match(vasim_50_w_match_126) ,
                .active_state(vasim_50_w_out_126));




/*wire vasim_50_w_out_127;
*/

wire vasim_50_lut_match_127;
wire vasim_50_w_match_127;

    
    
    

LUT_Match_vasim_50_127 #(8) lut_match_vasim_50_127(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_127));


assign vasim_50_w_match_127 = vasim_50_lut_match_127 ;

STE #(.fan_in(1)) vasim_50_ste_127 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_126 }),
                .match(vasim_50_w_match_127) ,
                .active_state(vasim_50_w_out_127));




/*wire vasim_50_w_out_128;
*/

wire vasim_50_lut_match_128;
wire vasim_50_w_match_128;

    
    
    

LUT_Match_vasim_50_128 #(8) lut_match_vasim_50_128(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_128));


assign vasim_50_w_match_128 = vasim_50_lut_match_128 ;

STE #(.fan_in(1)) vasim_50_ste_128 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_127 }),
                .match(vasim_50_w_match_128) ,
                .active_state(vasim_50_w_out_128));




/*wire vasim_50_w_out_129;
*/

wire vasim_50_lut_match_129;
wire vasim_50_w_match_129;

    
    
    

LUT_Match_vasim_50_129 #(8) lut_match_vasim_50_129(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_129));


assign vasim_50_w_match_129 = vasim_50_lut_match_129 ;

STE #(.fan_in(1)) vasim_50_ste_129 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_128 }),
                .match(vasim_50_w_match_129) ,
                .active_state(vasim_50_w_out_129));




/*wire vasim_50_w_out_130;
*/

wire vasim_50_lut_match_130;
wire vasim_50_w_match_130;

    
    
    

LUT_Match_vasim_50_130 #(8) lut_match_vasim_50_130(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_130));


assign vasim_50_w_match_130 = vasim_50_lut_match_130 ;

STE #(.fan_in(1)) vasim_50_ste_130 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_129 }),
                .match(vasim_50_w_match_130) ,
                .active_state(vasim_50_w_out_130));




/*wire vasim_50_w_out_131;
*/

wire vasim_50_lut_match_131;
wire vasim_50_w_match_131;

    
    
    

LUT_Match_vasim_50_131 #(8) lut_match_vasim_50_131(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_131));


assign vasim_50_w_match_131 = vasim_50_lut_match_131 ;

STE #(.fan_in(1)) vasim_50_ste_131 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_130 }),
                .match(vasim_50_w_match_131) ,
                .active_state(vasim_50_w_out_131));




/*wire vasim_50_w_out_132;
*/

wire vasim_50_lut_match_132;
wire vasim_50_w_match_132;

    
    
    

LUT_Match_vasim_50_132 #(8) lut_match_vasim_50_132(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_132));


assign vasim_50_w_match_132 = vasim_50_lut_match_132 ;

STE #(.fan_in(1)) vasim_50_ste_132 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_131 }),
                .match(vasim_50_w_match_132) ,
                .active_state(vasim_50_w_out_132));




/*wire vasim_50_w_out_133;
*/

wire vasim_50_lut_match_133;
wire vasim_50_w_match_133;

    
    
    

LUT_Match_vasim_50_133 #(8) lut_match_vasim_50_133(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_133));


assign vasim_50_w_match_133 = vasim_50_lut_match_133 ;

STE #(.fan_in(1)) vasim_50_ste_133 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_122 }),
                .match(vasim_50_w_match_133) ,
                .active_state(vasim_50_w_out_133));




/*wire vasim_50_w_out_134;
*/

wire vasim_50_lut_match_134;
wire vasim_50_w_match_134;

    
    
    

LUT_Match_vasim_50_134 #(8) lut_match_vasim_50_134(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_134));


assign vasim_50_w_match_134 = vasim_50_lut_match_134 ;

STE #(.fan_in(1)) vasim_50_ste_134 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_132 }),
                .match(vasim_50_w_match_134) ,
                .active_state(vasim_50_w_out_134));




/*wire vasim_50_w_out_135;
*/

wire vasim_50_lut_match_135;
wire vasim_50_w_match_135;

    
    
    

LUT_Match_vasim_50_135 #(8) lut_match_vasim_50_135(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_135));


assign vasim_50_w_match_135 = vasim_50_lut_match_135 ;

STE #(.fan_in(1)) vasim_50_ste_135 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_134 }),
                .match(vasim_50_w_match_135) ,
                .active_state(vasim_50_w_out_135));




/*wire vasim_50_w_out_136;
*/

wire vasim_50_lut_match_136;
wire vasim_50_w_match_136;

    
    
    

LUT_Match_vasim_50_136 #(8) lut_match_vasim_50_136(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_136));


assign vasim_50_w_match_136 = vasim_50_lut_match_136 ;

STE #(.fan_in(1)) vasim_50_ste_136 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_135 }),
                .match(vasim_50_w_match_136) ,
                .active_state(vasim_50_w_out_136));




/*wire vasim_50_w_out_137;
*/

wire vasim_50_lut_match_137;
wire vasim_50_w_match_137;

    
    
    

LUT_Match_vasim_50_137 #(8) lut_match_vasim_50_137(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_137));


assign vasim_50_w_match_137 = vasim_50_lut_match_137 ;

STE #(.fan_in(1)) vasim_50_ste_137 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_136 }),
                .match(vasim_50_w_match_137) ,
                .active_state(vasim_50_w_out_137));




/*wire vasim_50_w_out_138;
*/

wire vasim_50_lut_match_138;
wire vasim_50_w_match_138;

    
    
    

LUT_Match_vasim_50_138 #(8) lut_match_vasim_50_138(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_138));


assign vasim_50_w_match_138 = vasim_50_lut_match_138 ;

STE #(.fan_in(1)) vasim_50_ste_138 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_137 }),
                .match(vasim_50_w_match_138) ,
                .active_state(vasim_50_w_out_138));




/*wire vasim_50_w_out_139;
*/

wire vasim_50_lut_match_139;
wire vasim_50_w_match_139;

    
    
    

LUT_Match_vasim_50_139 #(8) lut_match_vasim_50_139(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_139));


assign vasim_50_w_match_139 = vasim_50_lut_match_139 ;

STE #(.fan_in(1)) vasim_50_ste_139 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_138 }),
                .match(vasim_50_w_match_139) ,
                .active_state(vasim_50_w_out_139));




/*wire vasim_50_w_out_140;
*/

wire vasim_50_lut_match_140;
wire vasim_50_w_match_140;

    
    
    

LUT_Match_vasim_50_140 #(8) lut_match_vasim_50_140(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_140));


assign vasim_50_w_match_140 = vasim_50_lut_match_140 ;

STE #(.fan_in(1)) vasim_50_ste_140 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_139 }),
                .match(vasim_50_w_match_140) ,
                .active_state(vasim_50_w_out_140));




/*wire vasim_50_w_out_141;
*/

wire vasim_50_lut_match_141;
wire vasim_50_w_match_141;

    
    
    

LUT_Match_vasim_50_141 #(8) lut_match_vasim_50_141(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_141));


assign vasim_50_w_match_141 = vasim_50_lut_match_141 ;

STE #(.fan_in(1)) vasim_50_ste_141 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_140 }),
                .match(vasim_50_w_match_141) ,
                .active_state(vasim_50_w_out_141));




/*wire vasim_50_w_out_142;
*/

wire vasim_50_lut_match_142;
wire vasim_50_w_match_142;

    
    
    

LUT_Match_vasim_50_142 #(8) lut_match_vasim_50_142(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_142));


assign vasim_50_w_match_142 = vasim_50_lut_match_142 ;

STE #(.fan_in(1)) vasim_50_ste_142 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_141 }),
                .match(vasim_50_w_match_142) ,
                .active_state(vasim_50_w_out_142));




/*wire vasim_50_w_out_143;
*/

wire vasim_50_lut_match_143;
wire vasim_50_w_match_143;

    
    
    

LUT_Match_vasim_50_143 #(8) lut_match_vasim_50_143(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_143));


assign vasim_50_w_match_143 = vasim_50_lut_match_143 ;

STE #(.fan_in(1)) vasim_50_ste_143 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_142 }),
                .match(vasim_50_w_match_143) ,
                .active_state(vasim_50_w_out_143));




/*wire vasim_50_w_out_144;
*/

wire vasim_50_lut_match_144;
wire vasim_50_w_match_144;

    
    
    

LUT_Match_vasim_50_144 #(8) lut_match_vasim_50_144(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_144));


assign vasim_50_w_match_144 = vasim_50_lut_match_144 ;

STE #(.fan_in(1)) vasim_50_ste_144 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_133 }),
                .match(vasim_50_w_match_144) ,
                .active_state(vasim_50_w_out_144));




/*wire vasim_50_w_out_145;
*/

wire vasim_50_lut_match_145;
wire vasim_50_w_match_145;

    
    
    

LUT_Match_vasim_50_145 #(8) lut_match_vasim_50_145(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_145));


assign vasim_50_w_match_145 = vasim_50_lut_match_145 ;

STE #(.fan_in(1)) vasim_50_ste_145 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_143 }),
                .match(vasim_50_w_match_145) ,
                .active_state(vasim_50_w_out_145));




/*wire vasim_50_w_out_146;
*/

wire vasim_50_lut_match_146;
wire vasim_50_w_match_146;

    
    
    

LUT_Match_vasim_50_146 #(8) lut_match_vasim_50_146(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_146));


assign vasim_50_w_match_146 = vasim_50_lut_match_146 ;

STE #(.fan_in(1)) vasim_50_ste_146 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_145 }),
                .match(vasim_50_w_match_146) ,
                .active_state(vasim_50_w_out_146));




/*wire vasim_50_w_out_147;
*/

wire vasim_50_lut_match_147;
wire vasim_50_w_match_147;

    
    
    

LUT_Match_vasim_50_147 #(8) lut_match_vasim_50_147(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_147));


assign vasim_50_w_match_147 = vasim_50_lut_match_147 ;

STE #(.fan_in(1)) vasim_50_ste_147 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_146 }),
                .match(vasim_50_w_match_147) ,
                .active_state(vasim_50_w_out_147));




/*wire vasim_50_w_out_148;
*/

wire vasim_50_lut_match_148;
wire vasim_50_w_match_148;

    
    
    

LUT_Match_vasim_50_148 #(8) lut_match_vasim_50_148(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_148));


assign vasim_50_w_match_148 = vasim_50_lut_match_148 ;

STE #(.fan_in(1)) vasim_50_ste_148 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_147 }),
                .match(vasim_50_w_match_148) ,
                .active_state(vasim_50_w_out_148));




/*wire vasim_50_w_out_149;
*/

wire vasim_50_lut_match_149;
wire vasim_50_w_match_149;

    
    
    

LUT_Match_vasim_50_149 #(8) lut_match_vasim_50_149(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_149));


assign vasim_50_w_match_149 = vasim_50_lut_match_149 ;

STE #(.fan_in(1)) vasim_50_ste_149 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_148 }),
                .match(vasim_50_w_match_149) ,
                .active_state(vasim_50_w_out_149));




/*wire vasim_50_w_out_150;
*/

wire vasim_50_lut_match_150;
wire vasim_50_w_match_150;

    
    
    

LUT_Match_vasim_50_150 #(8) lut_match_vasim_50_150(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_150));


assign vasim_50_w_match_150 = vasim_50_lut_match_150 ;

STE #(.fan_in(1)) vasim_50_ste_150 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_149 }),
                .match(vasim_50_w_match_150) ,
                .active_state(vasim_50_w_out_150));




/*wire vasim_50_w_out_151;
*/

wire vasim_50_lut_match_151;
wire vasim_50_w_match_151;

    
    
    

LUT_Match_vasim_50_151 #(8) lut_match_vasim_50_151(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_151));


assign vasim_50_w_match_151 = vasim_50_lut_match_151 ;

STE #(.fan_in(1)) vasim_50_ste_151 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_150 }),
                .match(vasim_50_w_match_151) ,
                .active_state(vasim_50_w_out_151));




/*wire vasim_50_w_out_152;
*/

wire vasim_50_lut_match_152;
wire vasim_50_w_match_152;

    
    
    

LUT_Match_vasim_50_152 #(8) lut_match_vasim_50_152(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_152));


assign vasim_50_w_match_152 = vasim_50_lut_match_152 ;

STE #(.fan_in(1)) vasim_50_ste_152 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_151 }),
                .match(vasim_50_w_match_152) ,
                .active_state(vasim_50_w_out_152));




/*wire vasim_50_w_out_153;
*/

wire vasim_50_lut_match_153;
wire vasim_50_w_match_153;

    
    
    

LUT_Match_vasim_50_153 #(8) lut_match_vasim_50_153(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_153));


assign vasim_50_w_match_153 = vasim_50_lut_match_153 ;

STE #(.fan_in(1)) vasim_50_ste_153 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_152 }),
                .match(vasim_50_w_match_153) ,
                .active_state(vasim_50_w_out_153));




/*wire vasim_50_w_out_154;
*/

wire vasim_50_lut_match_154;
wire vasim_50_w_match_154;

    
    
    

LUT_Match_vasim_50_154 #(8) lut_match_vasim_50_154(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_154));


assign vasim_50_w_match_154 = vasim_50_lut_match_154 ;

STE #(.fan_in(1)) vasim_50_ste_154 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_153 }),
                .match(vasim_50_w_match_154) ,
                .active_state(vasim_50_w_out_154));




/*wire vasim_50_w_out_155;
*/

wire vasim_50_lut_match_155;
wire vasim_50_w_match_155;

    
    
    

LUT_Match_vasim_50_155 #(8) lut_match_vasim_50_155(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_155));


assign vasim_50_w_match_155 = vasim_50_lut_match_155 ;

STE #(.fan_in(1)) vasim_50_ste_155 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_144 }),
                .match(vasim_50_w_match_155) ,
                .active_state(vasim_50_w_out_155));




/*wire vasim_50_w_out_156;
*/

wire vasim_50_lut_match_156;
wire vasim_50_w_match_156;

    
    
    

LUT_Match_vasim_50_156 #(8) lut_match_vasim_50_156(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_156));


assign vasim_50_w_match_156 = vasim_50_lut_match_156 ;

STE #(.fan_in(1)) vasim_50_ste_156 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_154 }),
                .match(vasim_50_w_match_156) ,
                .active_state(vasim_50_w_out_156));




/*wire vasim_50_w_out_157;
*/

wire vasim_50_lut_match_157;
wire vasim_50_w_match_157;

    
    
    

LUT_Match_vasim_50_157 #(8) lut_match_vasim_50_157(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_157));


assign vasim_50_w_match_157 = vasim_50_lut_match_157 ;

STE #(.fan_in(1)) vasim_50_ste_157 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_156 }),
                .match(vasim_50_w_match_157) ,
                .active_state(vasim_50_w_out_157));




/*wire vasim_50_w_out_158;
*/

wire vasim_50_lut_match_158;
wire vasim_50_w_match_158;

    
    
    

LUT_Match_vasim_50_158 #(8) lut_match_vasim_50_158(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_158));


assign vasim_50_w_match_158 = vasim_50_lut_match_158 ;

STE #(.fan_in(1)) vasim_50_ste_158 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_157 }),
                .match(vasim_50_w_match_158) ,
                .active_state(vasim_50_w_out_158));




/*wire vasim_50_w_out_159;
*/

wire vasim_50_lut_match_159;
wire vasim_50_w_match_159;

    
    
    

LUT_Match_vasim_50_159 #(8) lut_match_vasim_50_159(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_159));


assign vasim_50_w_match_159 = vasim_50_lut_match_159 ;

STE #(.fan_in(1)) vasim_50_ste_159 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_158 }),
                .match(vasim_50_w_match_159) ,
                .active_state(vasim_50_w_out_159));




/*wire vasim_50_w_out_160;
*/

wire vasim_50_lut_match_160;
wire vasim_50_w_match_160;

    
    
    

LUT_Match_vasim_50_160 #(8) lut_match_vasim_50_160(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_160));


assign vasim_50_w_match_160 = vasim_50_lut_match_160 ;

STE #(.fan_in(1)) vasim_50_ste_160 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_159 }),
                .match(vasim_50_w_match_160) ,
                .active_state(vasim_50_w_out_160));




/*wire vasim_50_w_out_161;
*/

wire vasim_50_lut_match_161;
wire vasim_50_w_match_161;

    
    
    

LUT_Match_vasim_50_161 #(8) lut_match_vasim_50_161(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_161));


assign vasim_50_w_match_161 = vasim_50_lut_match_161 ;

STE #(.fan_in(1)) vasim_50_ste_161 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_160 }),
                .match(vasim_50_w_match_161) ,
                .active_state(vasim_50_w_out_161));




/*wire vasim_50_w_out_162;
*/

wire vasim_50_lut_match_162;
wire vasim_50_w_match_162;

    
    
    

LUT_Match_vasim_50_162 #(8) lut_match_vasim_50_162(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_162));


assign vasim_50_w_match_162 = vasim_50_lut_match_162 ;

STE #(.fan_in(1)) vasim_50_ste_162 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_161 }),
                .match(vasim_50_w_match_162) ,
                .active_state(vasim_50_w_out_162));




/*wire vasim_50_w_out_163;
*/

wire vasim_50_lut_match_163;
wire vasim_50_w_match_163;

    
    
    

LUT_Match_vasim_50_163 #(8) lut_match_vasim_50_163(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_163));


assign vasim_50_w_match_163 = vasim_50_lut_match_163 ;

STE #(.fan_in(1)) vasim_50_ste_163 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_162 }),
                .match(vasim_50_w_match_163) ,
                .active_state(vasim_50_w_out_163));




/*wire vasim_50_w_out_164;
*/

wire vasim_50_lut_match_164;
wire vasim_50_w_match_164;

    
    
    

LUT_Match_vasim_50_164 #(8) lut_match_vasim_50_164(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_164));


assign vasim_50_w_match_164 = vasim_50_lut_match_164 ;

STE #(.fan_in(1)) vasim_50_ste_164 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_163 }),
                .match(vasim_50_w_match_164) ,
                .active_state(vasim_50_w_out_164));




/*wire vasim_50_w_out_165;
*/

wire vasim_50_lut_match_165;
wire vasim_50_w_match_165;

    
    
    

LUT_Match_vasim_50_165 #(8) lut_match_vasim_50_165(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_165));


assign vasim_50_w_match_165 = vasim_50_lut_match_165 ;

STE #(.fan_in(1)) vasim_50_ste_165 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_164 }),
                .match(vasim_50_w_match_165) ,
                .active_state(vasim_50_w_out_165));




/*wire vasim_50_w_out_166;
*/

wire vasim_50_lut_match_166;
wire vasim_50_w_match_166;

    
    
    

LUT_Match_vasim_50_166 #(8) lut_match_vasim_50_166(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_166));


assign vasim_50_w_match_166 = vasim_50_lut_match_166 ;

STE #(.fan_in(1)) vasim_50_ste_166 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_155 }),
                .match(vasim_50_w_match_166) ,
                .active_state(vasim_50_w_out_166));




/*wire vasim_50_w_out_167;
*/

wire vasim_50_lut_match_167;
wire vasim_50_w_match_167;

    
    
    

LUT_Match_vasim_50_167 #(8) lut_match_vasim_50_167(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_167));


assign vasim_50_w_match_167 = vasim_50_lut_match_167 ;

STE #(.fan_in(1)) vasim_50_ste_167 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_165 }),
                .match(vasim_50_w_match_167) ,
                .active_state(vasim_50_w_out_167));




/*wire vasim_50_w_out_168;
*/

wire vasim_50_lut_match_168;
wire vasim_50_w_match_168;

    
    
    

LUT_Match_vasim_50_168 #(8) lut_match_vasim_50_168(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_168));


assign vasim_50_w_match_168 = vasim_50_lut_match_168 ;

STE #(.fan_in(1)) vasim_50_ste_168 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_167 }),
                .match(vasim_50_w_match_168) ,
                .active_state(vasim_50_w_out_168));




/*wire vasim_50_w_out_169;
*/

wire vasim_50_lut_match_169;
wire vasim_50_w_match_169;

    
    
    

LUT_Match_vasim_50_169 #(8) lut_match_vasim_50_169(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_169));


assign vasim_50_w_match_169 = vasim_50_lut_match_169 ;

STE #(.fan_in(1)) vasim_50_ste_169 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_168 }),
                .match(vasim_50_w_match_169) ,
                .active_state(vasim_50_w_out_169));




/*wire vasim_50_w_out_170;
*/

wire vasim_50_lut_match_170;
wire vasim_50_w_match_170;

    
    
    

LUT_Match_vasim_50_170 #(8) lut_match_vasim_50_170(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_170));


assign vasim_50_w_match_170 = vasim_50_lut_match_170 ;

STE #(.fan_in(1)) vasim_50_ste_170 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_169 }),
                .match(vasim_50_w_match_170) ,
                .active_state(vasim_50_w_out_170));




/*wire vasim_50_w_out_171;
*/

wire vasim_50_lut_match_171;
wire vasim_50_w_match_171;

    
    
    

LUT_Match_vasim_50_171 #(8) lut_match_vasim_50_171(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_171));


assign vasim_50_w_match_171 = vasim_50_lut_match_171 ;

STE #(.fan_in(1)) vasim_50_ste_171 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_170 }),
                .match(vasim_50_w_match_171) ,
                .active_state(vasim_50_w_out_171));




/*wire vasim_50_w_out_172;
*/

wire vasim_50_lut_match_172;
wire vasim_50_w_match_172;

    
    
    

LUT_Match_vasim_50_172 #(8) lut_match_vasim_50_172(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_172));


assign vasim_50_w_match_172 = vasim_50_lut_match_172 ;

STE #(.fan_in(1)) vasim_50_ste_172 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_171 }),
                .match(vasim_50_w_match_172) ,
                .active_state(vasim_50_w_out_172));




/*wire vasim_50_w_out_173;
*/

wire vasim_50_lut_match_173;
wire vasim_50_w_match_173;

    
    
    

LUT_Match_vasim_50_173 #(8) lut_match_vasim_50_173(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_173));


assign vasim_50_w_match_173 = vasim_50_lut_match_173 ;

STE #(.fan_in(1)) vasim_50_ste_173 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_172 }),
                .match(vasim_50_w_match_173) ,
                .active_state(vasim_50_w_out_173));




/*wire vasim_50_w_out_174;
*/

wire vasim_50_lut_match_174;
wire vasim_50_w_match_174;

    
    
    

LUT_Match_vasim_50_174 #(8) lut_match_vasim_50_174(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_174));


assign vasim_50_w_match_174 = vasim_50_lut_match_174 ;

STE #(.fan_in(2)) vasim_50_ste_174 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_173, vasim_50_w_out_174 }),
                .match(vasim_50_w_match_174) ,
                .active_state(vasim_50_w_out_174));




/*wire vasim_50_w_out_175;
*/

wire vasim_50_lut_match_175;
wire vasim_50_w_match_175;

    
    
    

LUT_Match_vasim_50_175 #(8) lut_match_vasim_50_175(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_175));


assign vasim_50_w_match_175 = vasim_50_lut_match_175 ;

STE #(.fan_in(1)) vasim_50_ste_175 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_174 }),
                .match(vasim_50_w_match_175) ,
                .active_state(vasim_50_w_out_175));




/*wire vasim_50_w_out_176;
*/

wire vasim_50_lut_match_176;
wire vasim_50_w_match_176;

    
    
    

LUT_Match_vasim_50_176 #(8) lut_match_vasim_50_176(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_176));


assign vasim_50_w_match_176 = vasim_50_lut_match_176 ;

STE #(.fan_in(1)) vasim_50_ste_176 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_175 }),
                .match(vasim_50_w_match_176) ,
                .active_state(vasim_50_w_out_176));




/*wire vasim_50_w_out_177;
*/

wire vasim_50_lut_match_177;
wire vasim_50_w_match_177;

    
    
    

LUT_Match_vasim_50_177 #(8) lut_match_vasim_50_177(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_177));


assign vasim_50_w_match_177 = vasim_50_lut_match_177 ;

STE #(.fan_in(1)) vasim_50_ste_177 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_166 }),
                .match(vasim_50_w_match_177) ,
                .active_state(vasim_50_w_out_177));




/*wire vasim_50_w_out_178;
*/

wire vasim_50_lut_match_178;
wire vasim_50_w_match_178;

    
    
    

LUT_Match_vasim_50_178 #(8) lut_match_vasim_50_178(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_178));


assign vasim_50_w_match_178 = vasim_50_lut_match_178 ;

STE #(.fan_in(1)) vasim_50_ste_178 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_176 }),
                .match(vasim_50_w_match_178) ,
                .active_state(vasim_50_w_out_178));




/**/

wire vasim_50_lut_match_179;
wire vasim_50_w_match_179;

    
    
    

LUT_Match_vasim_50_179 #(8) lut_match_vasim_50_179(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_179));


assign vasim_50_w_match_179 = vasim_50_lut_match_179 ;

STE #(.fan_in(1)) vasim_50_ste_179 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_178 }),
                .match(vasim_50_w_match_179) ,
                .active_state(vasim_50_w_out_179));




/*wire vasim_50_w_out_180;
*/

wire vasim_50_lut_match_180;
wire vasim_50_w_match_180;

    
    
    

LUT_Match_vasim_50_180 #(8) lut_match_vasim_50_180(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_180));


assign vasim_50_w_match_180 = vasim_50_lut_match_180 ;

STE #(.fan_in(1)) vasim_50_ste_180 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_177 }),
                .match(vasim_50_w_match_180) ,
                .active_state(vasim_50_w_out_180));




/*wire vasim_50_w_out_181;
*/

wire vasim_50_lut_match_181;
wire vasim_50_w_match_181;

    
    
    

LUT_Match_vasim_50_181 #(8) lut_match_vasim_50_181(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_181));


assign vasim_50_w_match_181 = vasim_50_lut_match_181 ;

STE #(.fan_in(1)) vasim_50_ste_181 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_180 }),
                .match(vasim_50_w_match_181) ,
                .active_state(vasim_50_w_out_181));




/*wire vasim_50_w_out_182;
*/

wire vasim_50_lut_match_182;
wire vasim_50_w_match_182;

    
    
    

LUT_Match_vasim_50_182 #(8) lut_match_vasim_50_182(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_182));


assign vasim_50_w_match_182 = vasim_50_lut_match_182 ;

STE #(.fan_in(1)) vasim_50_ste_182 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_181 }),
                .match(vasim_50_w_match_182) ,
                .active_state(vasim_50_w_out_182));




/*wire vasim_50_w_out_183;
*/

wire vasim_50_lut_match_183;
wire vasim_50_w_match_183;

    
    
    

LUT_Match_vasim_50_183 #(8) lut_match_vasim_50_183(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_183));


assign vasim_50_w_match_183 = vasim_50_lut_match_183 ;

STE #(.fan_in(1)) vasim_50_ste_183 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_182 }),
                .match(vasim_50_w_match_183) ,
                .active_state(vasim_50_w_out_183));




/*wire vasim_50_w_out_184;
*/

wire vasim_50_lut_match_184;
wire vasim_50_w_match_184;

    
    
    

LUT_Match_vasim_50_184 #(8) lut_match_vasim_50_184(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_184));


assign vasim_50_w_match_184 = vasim_50_lut_match_184 ;

STE #(.fan_in(1)) vasim_50_ste_184 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_183 }),
                .match(vasim_50_w_match_184) ,
                .active_state(vasim_50_w_out_184));




/*wire vasim_50_w_out_185;
*/

wire vasim_50_lut_match_185;
wire vasim_50_w_match_185;

    
    
    

LUT_Match_vasim_50_185 #(8) lut_match_vasim_50_185(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_185));


assign vasim_50_w_match_185 = vasim_50_lut_match_185 ;

STE #(.fan_in(1)) vasim_50_ste_185 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_184 }),
                .match(vasim_50_w_match_185) ,
                .active_state(vasim_50_w_out_185));




/*wire vasim_50_w_out_186;
*/

wire vasim_50_lut_match_186;
wire vasim_50_w_match_186;

    
    
    

LUT_Match_vasim_50_186 #(8) lut_match_vasim_50_186(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_186));


assign vasim_50_w_match_186 = vasim_50_lut_match_186 ;

STE #(.fan_in(1)) vasim_50_ste_186 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_185 }),
                .match(vasim_50_w_match_186) ,
                .active_state(vasim_50_w_out_186));




/*wire vasim_50_w_out_187;
*/

wire vasim_50_lut_match_187;
wire vasim_50_w_match_187;

    
    
    

LUT_Match_vasim_50_187 #(8) lut_match_vasim_50_187(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_187));


assign vasim_50_w_match_187 = vasim_50_lut_match_187 ;

STE #(.fan_in(1)) vasim_50_ste_187 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_186 }),
                .match(vasim_50_w_match_187) ,
                .active_state(vasim_50_w_out_187));




/*wire vasim_50_w_out_188;
*/

wire vasim_50_lut_match_188;
wire vasim_50_w_match_188;

    
    
    

LUT_Match_vasim_50_188 #(8) lut_match_vasim_50_188(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_188));


assign vasim_50_w_match_188 = vasim_50_lut_match_188 ;

STE #(.fan_in(1)) vasim_50_ste_188 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_187 }),
                .match(vasim_50_w_match_188) ,
                .active_state(vasim_50_w_out_188));




/*wire vasim_50_w_out_189;
*/

wire vasim_50_lut_match_189;
wire vasim_50_w_match_189;

    
    
    

LUT_Match_vasim_50_189 #(8) lut_match_vasim_50_189(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_189));


assign vasim_50_w_match_189 = vasim_50_lut_match_189 ;

STE #(.fan_in(1)) vasim_50_ste_189 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_188 }),
                .match(vasim_50_w_match_189) ,
                .active_state(vasim_50_w_out_189));




/*wire vasim_50_w_out_190;
*/

wire vasim_50_lut_match_190;
wire vasim_50_w_match_190;

    
    
    

LUT_Match_vasim_50_190 #(8) lut_match_vasim_50_190(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_190));


assign vasim_50_w_match_190 = vasim_50_lut_match_190 ;

STE #(.fan_in(1)) vasim_50_ste_190 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_189 }),
                .match(vasim_50_w_match_190) ,
                .active_state(vasim_50_w_out_190));




/*wire vasim_50_w_out_191;
*/

wire vasim_50_lut_match_191;
wire vasim_50_w_match_191;

    
    
    

LUT_Match_vasim_50_191 #(8) lut_match_vasim_50_191(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_191));


assign vasim_50_w_match_191 = vasim_50_lut_match_191 ;

STE #(.fan_in(1)) vasim_50_ste_191 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_190 }),
                .match(vasim_50_w_match_191) ,
                .active_state(vasim_50_w_out_191));




/*wire vasim_50_w_out_192;
*/

wire vasim_50_lut_match_192;
wire vasim_50_w_match_192;

    
    
    

LUT_Match_vasim_50_192 #(8) lut_match_vasim_50_192(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_192));


assign vasim_50_w_match_192 = vasim_50_lut_match_192 ;

STE #(.fan_in(1)) vasim_50_ste_192 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_191 }),
                .match(vasim_50_w_match_192) ,
                .active_state(vasim_50_w_out_192));




/*wire vasim_50_w_out_193;
*/

wire vasim_50_lut_match_193;
wire vasim_50_w_match_193;

    
    
    
            

LUT_Match_vasim_50_193 #(8) lut_match_vasim_50_193(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_193));


assign vasim_50_w_match_193 = vasim_50_lut_match_193 ;

STE #(.fan_in(1),.START_TYPE(2)) vasim_50_ste_193 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ all_input }),
                .match(vasim_50_w_match_193) ,
                .active_state(vasim_50_w_out_193));




/*wire vasim_50_w_out_194;
*/

wire vasim_50_lut_match_194;
wire vasim_50_w_match_194;

    
    
    

LUT_Match_vasim_50_194 #(8) lut_match_vasim_50_194(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_194));


assign vasim_50_w_match_194 = vasim_50_lut_match_194 ;

STE #(.fan_in(1)) vasim_50_ste_194 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_192 }),
                .match(vasim_50_w_match_194) ,
                .active_state(vasim_50_w_out_194));




/*wire vasim_50_w_out_195;
*/

wire vasim_50_lut_match_195;
wire vasim_50_w_match_195;

    
    
    

LUT_Match_vasim_50_195 #(8) lut_match_vasim_50_195(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_195));


assign vasim_50_w_match_195 = vasim_50_lut_match_195 ;

STE #(.fan_in(1)) vasim_50_ste_195 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_194 }),
                .match(vasim_50_w_match_195) ,
                .active_state(vasim_50_w_out_195));




/*wire vasim_50_w_out_196;
*/

wire vasim_50_lut_match_196;
wire vasim_50_w_match_196;

    
    
    

LUT_Match_vasim_50_196 #(8) lut_match_vasim_50_196(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_196));


assign vasim_50_w_match_196 = vasim_50_lut_match_196 ;

STE #(.fan_in(1)) vasim_50_ste_196 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_195 }),
                .match(vasim_50_w_match_196) ,
                .active_state(vasim_50_w_out_196));




/*wire vasim_50_w_out_197;
*/

wire vasim_50_lut_match_197;
wire vasim_50_w_match_197;

    
    
    

LUT_Match_vasim_50_197 #(8) lut_match_vasim_50_197(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_197));


assign vasim_50_w_match_197 = vasim_50_lut_match_197 ;

STE #(.fan_in(1)) vasim_50_ste_197 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_196 }),
                .match(vasim_50_w_match_197) ,
                .active_state(vasim_50_w_out_197));




/*wire vasim_50_w_out_198;
*/

wire vasim_50_lut_match_198;
wire vasim_50_w_match_198;

    
    
    

LUT_Match_vasim_50_198 #(8) lut_match_vasim_50_198(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_198));


assign vasim_50_w_match_198 = vasim_50_lut_match_198 ;

STE #(.fan_in(1)) vasim_50_ste_198 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_197 }),
                .match(vasim_50_w_match_198) ,
                .active_state(vasim_50_w_out_198));




/*wire vasim_50_w_out_199;
*/

wire vasim_50_lut_match_199;
wire vasim_50_w_match_199;

    
    
    

LUT_Match_vasim_50_199 #(8) lut_match_vasim_50_199(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_199));


assign vasim_50_w_match_199 = vasim_50_lut_match_199 ;

STE #(.fan_in(1)) vasim_50_ste_199 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_198 }),
                .match(vasim_50_w_match_199) ,
                .active_state(vasim_50_w_out_199));




/*wire vasim_50_w_out_200;
*/

wire vasim_50_lut_match_200;
wire vasim_50_w_match_200;

    
    
    

LUT_Match_vasim_50_200 #(8) lut_match_vasim_50_200(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_200));


assign vasim_50_w_match_200 = vasim_50_lut_match_200 ;

STE #(.fan_in(1)) vasim_50_ste_200 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_199 }),
                .match(vasim_50_w_match_200) ,
                .active_state(vasim_50_w_out_200));




/*wire vasim_50_w_out_201;
*/

wire vasim_50_lut_match_201;
wire vasim_50_w_match_201;

    
    
    

LUT_Match_vasim_50_201 #(8) lut_match_vasim_50_201(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_201));


assign vasim_50_w_match_201 = vasim_50_lut_match_201 ;

STE #(.fan_in(1)) vasim_50_ste_201 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_200 }),
                .match(vasim_50_w_match_201) ,
                .active_state(vasim_50_w_out_201));




/*wire vasim_50_w_out_202;
*/

wire vasim_50_lut_match_202;
wire vasim_50_w_match_202;

    
    
    

LUT_Match_vasim_50_202 #(8) lut_match_vasim_50_202(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_202));


assign vasim_50_w_match_202 = vasim_50_lut_match_202 ;

STE #(.fan_in(1)) vasim_50_ste_202 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_201 }),
                .match(vasim_50_w_match_202) ,
                .active_state(vasim_50_w_out_202));




/*wire vasim_50_w_out_203;
*/

wire vasim_50_lut_match_203;
wire vasim_50_w_match_203;

    
    
    

LUT_Match_vasim_50_203 #(8) lut_match_vasim_50_203(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_203));


assign vasim_50_w_match_203 = vasim_50_lut_match_203 ;

STE #(.fan_in(1)) vasim_50_ste_203 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_202 }),
                .match(vasim_50_w_match_203) ,
                .active_state(vasim_50_w_out_203));




/*wire vasim_50_w_out_204;
*/

wire vasim_50_lut_match_204;
wire vasim_50_w_match_204;

    
    
    

LUT_Match_vasim_50_204 #(8) lut_match_vasim_50_204(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_204));


assign vasim_50_w_match_204 = vasim_50_lut_match_204 ;

STE #(.fan_in(1)) vasim_50_ste_204 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_193 }),
                .match(vasim_50_w_match_204) ,
                .active_state(vasim_50_w_out_204));




/*wire vasim_50_w_out_205;
*/

wire vasim_50_lut_match_205;
wire vasim_50_w_match_205;

    
    
    

LUT_Match_vasim_50_205 #(8) lut_match_vasim_50_205(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_205));


assign vasim_50_w_match_205 = vasim_50_lut_match_205 ;

STE #(.fan_in(1)) vasim_50_ste_205 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_203 }),
                .match(vasim_50_w_match_205) ,
                .active_state(vasim_50_w_out_205));




/*wire vasim_50_w_out_206;
*/

wire vasim_50_lut_match_206;
wire vasim_50_w_match_206;

    
    
    

LUT_Match_vasim_50_206 #(8) lut_match_vasim_50_206(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_206));


assign vasim_50_w_match_206 = vasim_50_lut_match_206 ;

STE #(.fan_in(1)) vasim_50_ste_206 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_205 }),
                .match(vasim_50_w_match_206) ,
                .active_state(vasim_50_w_out_206));




/*wire vasim_50_w_out_207;
*/

wire vasim_50_lut_match_207;
wire vasim_50_w_match_207;

    
    
    

LUT_Match_vasim_50_207 #(8) lut_match_vasim_50_207(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_207));


assign vasim_50_w_match_207 = vasim_50_lut_match_207 ;

STE #(.fan_in(1)) vasim_50_ste_207 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_206 }),
                .match(vasim_50_w_match_207) ,
                .active_state(vasim_50_w_out_207));




/*wire vasim_50_w_out_208;
*/

wire vasim_50_lut_match_208;
wire vasim_50_w_match_208;

    
    
    

LUT_Match_vasim_50_208 #(8) lut_match_vasim_50_208(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_208));


assign vasim_50_w_match_208 = vasim_50_lut_match_208 ;

STE #(.fan_in(1)) vasim_50_ste_208 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_207 }),
                .match(vasim_50_w_match_208) ,
                .active_state(vasim_50_w_out_208));




/*wire vasim_50_w_out_209;
*/

wire vasim_50_lut_match_209;
wire vasim_50_w_match_209;

    
    
    

LUT_Match_vasim_50_209 #(8) lut_match_vasim_50_209(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_209));


assign vasim_50_w_match_209 = vasim_50_lut_match_209 ;

STE #(.fan_in(1)) vasim_50_ste_209 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_208 }),
                .match(vasim_50_w_match_209) ,
                .active_state(vasim_50_w_out_209));




/*wire vasim_50_w_out_210;
*/

wire vasim_50_lut_match_210;
wire vasim_50_w_match_210;

    
    
    

LUT_Match_vasim_50_210 #(8) lut_match_vasim_50_210(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_210));


assign vasim_50_w_match_210 = vasim_50_lut_match_210 ;

STE #(.fan_in(1)) vasim_50_ste_210 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_209 }),
                .match(vasim_50_w_match_210) ,
                .active_state(vasim_50_w_out_210));




/*wire vasim_50_w_out_211;
*/

wire vasim_50_lut_match_211;
wire vasim_50_w_match_211;

    
    
    

LUT_Match_vasim_50_211 #(8) lut_match_vasim_50_211(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_211));


assign vasim_50_w_match_211 = vasim_50_lut_match_211 ;

STE #(.fan_in(1)) vasim_50_ste_211 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_210 }),
                .match(vasim_50_w_match_211) ,
                .active_state(vasim_50_w_out_211));




/*wire vasim_50_w_out_212;
*/

wire vasim_50_lut_match_212;
wire vasim_50_w_match_212;

    
    
    

LUT_Match_vasim_50_212 #(8) lut_match_vasim_50_212(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_212));


assign vasim_50_w_match_212 = vasim_50_lut_match_212 ;

STE #(.fan_in(1)) vasim_50_ste_212 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_211 }),
                .match(vasim_50_w_match_212) ,
                .active_state(vasim_50_w_out_212));




/*wire vasim_50_w_out_213;
*/

wire vasim_50_lut_match_213;
wire vasim_50_w_match_213;

    
    
    

LUT_Match_vasim_50_213 #(8) lut_match_vasim_50_213(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_213));


assign vasim_50_w_match_213 = vasim_50_lut_match_213 ;

STE #(.fan_in(1)) vasim_50_ste_213 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_212 }),
                .match(vasim_50_w_match_213) ,
                .active_state(vasim_50_w_out_213));




/*wire vasim_50_w_out_214;
*/

wire vasim_50_lut_match_214;
wire vasim_50_w_match_214;

    
    
    

LUT_Match_vasim_50_214 #(8) lut_match_vasim_50_214(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_214));


assign vasim_50_w_match_214 = vasim_50_lut_match_214 ;

STE #(.fan_in(1)) vasim_50_ste_214 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_213 }),
                .match(vasim_50_w_match_214) ,
                .active_state(vasim_50_w_out_214));




/*wire vasim_50_w_out_215;
*/

wire vasim_50_lut_match_215;
wire vasim_50_w_match_215;

    
    
    

LUT_Match_vasim_50_215 #(8) lut_match_vasim_50_215(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_215));


assign vasim_50_w_match_215 = vasim_50_lut_match_215 ;

STE #(.fan_in(1)) vasim_50_ste_215 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_204 }),
                .match(vasim_50_w_match_215) ,
                .active_state(vasim_50_w_out_215));




/*wire vasim_50_w_out_216;
*/

wire vasim_50_lut_match_216;
wire vasim_50_w_match_216;

    
    
    

LUT_Match_vasim_50_216 #(8) lut_match_vasim_50_216(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_216));


assign vasim_50_w_match_216 = vasim_50_lut_match_216 ;

STE #(.fan_in(1)) vasim_50_ste_216 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_214 }),
                .match(vasim_50_w_match_216) ,
                .active_state(vasim_50_w_out_216));




/*wire vasim_50_w_out_217;
*/

wire vasim_50_lut_match_217;
wire vasim_50_w_match_217;

    
    
    

LUT_Match_vasim_50_217 #(8) lut_match_vasim_50_217(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_217));


assign vasim_50_w_match_217 = vasim_50_lut_match_217 ;

STE #(.fan_in(1)) vasim_50_ste_217 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_216 }),
                .match(vasim_50_w_match_217) ,
                .active_state(vasim_50_w_out_217));




/*wire vasim_50_w_out_218;
*/

wire vasim_50_lut_match_218;
wire vasim_50_w_match_218;

    
    
    

LUT_Match_vasim_50_218 #(8) lut_match_vasim_50_218(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_218));


assign vasim_50_w_match_218 = vasim_50_lut_match_218 ;

STE #(.fan_in(1)) vasim_50_ste_218 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_217 }),
                .match(vasim_50_w_match_218) ,
                .active_state(vasim_50_w_out_218));




/*wire vasim_50_w_out_219;
*/

wire vasim_50_lut_match_219;
wire vasim_50_w_match_219;

    
    
    

LUT_Match_vasim_50_219 #(8) lut_match_vasim_50_219(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_219));


assign vasim_50_w_match_219 = vasim_50_lut_match_219 ;

STE #(.fan_in(1)) vasim_50_ste_219 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_218 }),
                .match(vasim_50_w_match_219) ,
                .active_state(vasim_50_w_out_219));




/*wire vasim_50_w_out_220;
*/

wire vasim_50_lut_match_220;
wire vasim_50_w_match_220;

    
    
    

LUT_Match_vasim_50_220 #(8) lut_match_vasim_50_220(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_220));


assign vasim_50_w_match_220 = vasim_50_lut_match_220 ;

STE #(.fan_in(1)) vasim_50_ste_220 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_219 }),
                .match(vasim_50_w_match_220) ,
                .active_state(vasim_50_w_out_220));




/*wire vasim_50_w_out_221;
*/

wire vasim_50_lut_match_221;
wire vasim_50_w_match_221;

    
    
    

LUT_Match_vasim_50_221 #(8) lut_match_vasim_50_221(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_221));


assign vasim_50_w_match_221 = vasim_50_lut_match_221 ;

STE #(.fan_in(1)) vasim_50_ste_221 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_220 }),
                .match(vasim_50_w_match_221) ,
                .active_state(vasim_50_w_out_221));




/*wire vasim_50_w_out_222;
*/

wire vasim_50_lut_match_222;
wire vasim_50_w_match_222;

    
    
    

LUT_Match_vasim_50_222 #(8) lut_match_vasim_50_222(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_222));


assign vasim_50_w_match_222 = vasim_50_lut_match_222 ;

STE #(.fan_in(1)) vasim_50_ste_222 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_221 }),
                .match(vasim_50_w_match_222) ,
                .active_state(vasim_50_w_out_222));




/*wire vasim_50_w_out_223;
*/

wire vasim_50_lut_match_223;
wire vasim_50_w_match_223;

    
    
    

LUT_Match_vasim_50_223 #(8) lut_match_vasim_50_223(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_223));


assign vasim_50_w_match_223 = vasim_50_lut_match_223 ;

STE #(.fan_in(1)) vasim_50_ste_223 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_222 }),
                .match(vasim_50_w_match_223) ,
                .active_state(vasim_50_w_out_223));




/*wire vasim_50_w_out_224;
*/

wire vasim_50_lut_match_224;
wire vasim_50_w_match_224;

    
    
    

LUT_Match_vasim_50_224 #(8) lut_match_vasim_50_224(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_224));


assign vasim_50_w_match_224 = vasim_50_lut_match_224 ;

STE #(.fan_in(1)) vasim_50_ste_224 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_223 }),
                .match(vasim_50_w_match_224) ,
                .active_state(vasim_50_w_out_224));




/*wire vasim_50_w_out_225;
*/

wire vasim_50_lut_match_225;
wire vasim_50_w_match_225;

    
    
    

LUT_Match_vasim_50_225 #(8) lut_match_vasim_50_225(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_225));


assign vasim_50_w_match_225 = vasim_50_lut_match_225 ;

STE #(.fan_in(1)) vasim_50_ste_225 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_224 }),
                .match(vasim_50_w_match_225) ,
                .active_state(vasim_50_w_out_225));




/*wire vasim_50_w_out_226;
*/

wire vasim_50_lut_match_226;
wire vasim_50_w_match_226;

    
    
    

LUT_Match_vasim_50_226 #(8) lut_match_vasim_50_226(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_226));


assign vasim_50_w_match_226 = vasim_50_lut_match_226 ;

STE #(.fan_in(1)) vasim_50_ste_226 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_215 }),
                .match(vasim_50_w_match_226) ,
                .active_state(vasim_50_w_out_226));




/*wire vasim_50_w_out_227;
*/

wire vasim_50_lut_match_227;
wire vasim_50_w_match_227;

    
    
    

LUT_Match_vasim_50_227 #(8) lut_match_vasim_50_227(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_227));


assign vasim_50_w_match_227 = vasim_50_lut_match_227 ;

STE #(.fan_in(1)) vasim_50_ste_227 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_225 }),
                .match(vasim_50_w_match_227) ,
                .active_state(vasim_50_w_out_227));




/*wire vasim_50_w_out_228;
*/

wire vasim_50_lut_match_228;
wire vasim_50_w_match_228;

    
    
    

LUT_Match_vasim_50_228 #(8) lut_match_vasim_50_228(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_228));


assign vasim_50_w_match_228 = vasim_50_lut_match_228 ;

STE #(.fan_in(1)) vasim_50_ste_228 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_227 }),
                .match(vasim_50_w_match_228) ,
                .active_state(vasim_50_w_out_228));




/*wire vasim_50_w_out_229;
*/

wire vasim_50_lut_match_229;
wire vasim_50_w_match_229;

    
    
    

LUT_Match_vasim_50_229 #(8) lut_match_vasim_50_229(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_229));


assign vasim_50_w_match_229 = vasim_50_lut_match_229 ;

STE #(.fan_in(1)) vasim_50_ste_229 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_228 }),
                .match(vasim_50_w_match_229) ,
                .active_state(vasim_50_w_out_229));




/*wire vasim_50_w_out_230;
*/

wire vasim_50_lut_match_230;
wire vasim_50_w_match_230;

    
    
    

LUT_Match_vasim_50_230 #(8) lut_match_vasim_50_230(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_230));


assign vasim_50_w_match_230 = vasim_50_lut_match_230 ;

STE #(.fan_in(1)) vasim_50_ste_230 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_229 }),
                .match(vasim_50_w_match_230) ,
                .active_state(vasim_50_w_out_230));




/*wire vasim_50_w_out_231;
*/

wire vasim_50_lut_match_231;
wire vasim_50_w_match_231;

    
    
    

LUT_Match_vasim_50_231 #(8) lut_match_vasim_50_231(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_231));


assign vasim_50_w_match_231 = vasim_50_lut_match_231 ;

STE #(.fan_in(1)) vasim_50_ste_231 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_230 }),
                .match(vasim_50_w_match_231) ,
                .active_state(vasim_50_w_out_231));




/*wire vasim_50_w_out_232;
*/

wire vasim_50_lut_match_232;
wire vasim_50_w_match_232;

    
    
    

LUT_Match_vasim_50_232 #(8) lut_match_vasim_50_232(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_232));


assign vasim_50_w_match_232 = vasim_50_lut_match_232 ;

STE #(.fan_in(1)) vasim_50_ste_232 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_231 }),
                .match(vasim_50_w_match_232) ,
                .active_state(vasim_50_w_out_232));




/*wire vasim_50_w_out_233;
*/

wire vasim_50_lut_match_233;
wire vasim_50_w_match_233;

    
    
    

LUT_Match_vasim_50_233 #(8) lut_match_vasim_50_233(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_233));


assign vasim_50_w_match_233 = vasim_50_lut_match_233 ;

STE #(.fan_in(1)) vasim_50_ste_233 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_232 }),
                .match(vasim_50_w_match_233) ,
                .active_state(vasim_50_w_out_233));




/*wire vasim_50_w_out_234;
*/

wire vasim_50_lut_match_234;
wire vasim_50_w_match_234;

    
    
    

LUT_Match_vasim_50_234 #(8) lut_match_vasim_50_234(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_234));


assign vasim_50_w_match_234 = vasim_50_lut_match_234 ;

STE #(.fan_in(1)) vasim_50_ste_234 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_233 }),
                .match(vasim_50_w_match_234) ,
                .active_state(vasim_50_w_out_234));




/*wire vasim_50_w_out_235;
*/

wire vasim_50_lut_match_235;
wire vasim_50_w_match_235;

    
    
    

LUT_Match_vasim_50_235 #(8) lut_match_vasim_50_235(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_235));


assign vasim_50_w_match_235 = vasim_50_lut_match_235 ;

STE #(.fan_in(1)) vasim_50_ste_235 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_234 }),
                .match(vasim_50_w_match_235) ,
                .active_state(vasim_50_w_out_235));




/*wire vasim_50_w_out_236;
*/

wire vasim_50_lut_match_236;
wire vasim_50_w_match_236;

    
    
    

LUT_Match_vasim_50_236 #(8) lut_match_vasim_50_236(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_236));


assign vasim_50_w_match_236 = vasim_50_lut_match_236 ;

STE #(.fan_in(1)) vasim_50_ste_236 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_235 }),
                .match(vasim_50_w_match_236) ,
                .active_state(vasim_50_w_out_236));




/*wire vasim_50_w_out_237;
*/

wire vasim_50_lut_match_237;
wire vasim_50_w_match_237;

    
    
    

LUT_Match_vasim_50_237 #(8) lut_match_vasim_50_237(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_237));


assign vasim_50_w_match_237 = vasim_50_lut_match_237 ;

STE #(.fan_in(1)) vasim_50_ste_237 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_226 }),
                .match(vasim_50_w_match_237) ,
                .active_state(vasim_50_w_out_237));




/*wire vasim_50_w_out_238;
*/

wire vasim_50_lut_match_238;
wire vasim_50_w_match_238;

    
    
    

LUT_Match_vasim_50_238 #(8) lut_match_vasim_50_238(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_238));


assign vasim_50_w_match_238 = vasim_50_lut_match_238 ;

STE #(.fan_in(1)) vasim_50_ste_238 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_236 }),
                .match(vasim_50_w_match_238) ,
                .active_state(vasim_50_w_out_238));




/*wire vasim_50_w_out_239;
*/

wire vasim_50_lut_match_239;
wire vasim_50_w_match_239;

    
    
    

LUT_Match_vasim_50_239 #(8) lut_match_vasim_50_239(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_239));


assign vasim_50_w_match_239 = vasim_50_lut_match_239 ;

STE #(.fan_in(1)) vasim_50_ste_239 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_238 }),
                .match(vasim_50_w_match_239) ,
                .active_state(vasim_50_w_out_239));




/*wire vasim_50_w_out_240;
*/

wire vasim_50_lut_match_240;
wire vasim_50_w_match_240;

    
    
    

LUT_Match_vasim_50_240 #(8) lut_match_vasim_50_240(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_240));


assign vasim_50_w_match_240 = vasim_50_lut_match_240 ;

STE #(.fan_in(1)) vasim_50_ste_240 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_239 }),
                .match(vasim_50_w_match_240) ,
                .active_state(vasim_50_w_out_240));




/*wire vasim_50_w_out_241;
*/

wire vasim_50_lut_match_241;
wire vasim_50_w_match_241;

    
    
    

LUT_Match_vasim_50_241 #(8) lut_match_vasim_50_241(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_241));


assign vasim_50_w_match_241 = vasim_50_lut_match_241 ;

STE #(.fan_in(1)) vasim_50_ste_241 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_240 }),
                .match(vasim_50_w_match_241) ,
                .active_state(vasim_50_w_out_241));




/*wire vasim_50_w_out_242;
*/

wire vasim_50_lut_match_242;
wire vasim_50_w_match_242;

    
    
    

LUT_Match_vasim_50_242 #(8) lut_match_vasim_50_242(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_242));


assign vasim_50_w_match_242 = vasim_50_lut_match_242 ;

STE #(.fan_in(1)) vasim_50_ste_242 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_241 }),
                .match(vasim_50_w_match_242) ,
                .active_state(vasim_50_w_out_242));




/*wire vasim_50_w_out_243;
*/

wire vasim_50_lut_match_243;
wire vasim_50_w_match_243;

    
    
    

LUT_Match_vasim_50_243 #(8) lut_match_vasim_50_243(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_243));


assign vasim_50_w_match_243 = vasim_50_lut_match_243 ;

STE #(.fan_in(1)) vasim_50_ste_243 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_242 }),
                .match(vasim_50_w_match_243) ,
                .active_state(vasim_50_w_out_243));




/*wire vasim_50_w_out_244;
*/

wire vasim_50_lut_match_244;
wire vasim_50_w_match_244;

    
    
    

LUT_Match_vasim_50_244 #(8) lut_match_vasim_50_244(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_244));


assign vasim_50_w_match_244 = vasim_50_lut_match_244 ;

STE #(.fan_in(1)) vasim_50_ste_244 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_243 }),
                .match(vasim_50_w_match_244) ,
                .active_state(vasim_50_w_out_244));




/*wire vasim_50_w_out_245;
*/

wire vasim_50_lut_match_245;
wire vasim_50_w_match_245;

    
    
    

LUT_Match_vasim_50_245 #(8) lut_match_vasim_50_245(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_245));


assign vasim_50_w_match_245 = vasim_50_lut_match_245 ;

STE #(.fan_in(1)) vasim_50_ste_245 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_244 }),
                .match(vasim_50_w_match_245) ,
                .active_state(vasim_50_w_out_245));




/*wire vasim_50_w_out_246;
*/

wire vasim_50_lut_match_246;
wire vasim_50_w_match_246;

    
    
    

LUT_Match_vasim_50_246 #(8) lut_match_vasim_50_246(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_246));


assign vasim_50_w_match_246 = vasim_50_lut_match_246 ;

STE #(.fan_in(1)) vasim_50_ste_246 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_245 }),
                .match(vasim_50_w_match_246) ,
                .active_state(vasim_50_w_out_246));




/*wire vasim_50_w_out_247;
*/

wire vasim_50_lut_match_247;
wire vasim_50_w_match_247;

    
    
    

LUT_Match_vasim_50_247 #(8) lut_match_vasim_50_247(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_247));


assign vasim_50_w_match_247 = vasim_50_lut_match_247 ;

STE #(.fan_in(1)) vasim_50_ste_247 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_246 }),
                .match(vasim_50_w_match_247) ,
                .active_state(vasim_50_w_out_247));




/*wire vasim_50_w_out_248;
*/

wire vasim_50_lut_match_248;
wire vasim_50_w_match_248;

    
    
    

LUT_Match_vasim_50_248 #(8) lut_match_vasim_50_248(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_248));


assign vasim_50_w_match_248 = vasim_50_lut_match_248 ;

STE #(.fan_in(1)) vasim_50_ste_248 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_237 }),
                .match(vasim_50_w_match_248) ,
                .active_state(vasim_50_w_out_248));




/*wire vasim_50_w_out_249;
*/

wire vasim_50_lut_match_249;
wire vasim_50_w_match_249;

    
    
    

LUT_Match_vasim_50_249 #(8) lut_match_vasim_50_249(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_249));


assign vasim_50_w_match_249 = vasim_50_lut_match_249 ;

STE #(.fan_in(1)) vasim_50_ste_249 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_247 }),
                .match(vasim_50_w_match_249) ,
                .active_state(vasim_50_w_out_249));




/*wire vasim_50_w_out_250;
*/

wire vasim_50_lut_match_250;
wire vasim_50_w_match_250;

    
    
    

LUT_Match_vasim_50_250 #(8) lut_match_vasim_50_250(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_250));


assign vasim_50_w_match_250 = vasim_50_lut_match_250 ;

STE #(.fan_in(1)) vasim_50_ste_250 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_249 }),
                .match(vasim_50_w_match_250) ,
                .active_state(vasim_50_w_out_250));




/*wire vasim_50_w_out_251;
*/

wire vasim_50_lut_match_251;
wire vasim_50_w_match_251;

    
    
    

LUT_Match_vasim_50_251 #(8) lut_match_vasim_50_251(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_251));


assign vasim_50_w_match_251 = vasim_50_lut_match_251 ;

STE #(.fan_in(1)) vasim_50_ste_251 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_250 }),
                .match(vasim_50_w_match_251) ,
                .active_state(vasim_50_w_out_251));




/*wire vasim_50_w_out_252;
*/

wire vasim_50_lut_match_252;
wire vasim_50_w_match_252;

    
    
    

LUT_Match_vasim_50_252 #(8) lut_match_vasim_50_252(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_252));


assign vasim_50_w_match_252 = vasim_50_lut_match_252 ;

STE #(.fan_in(1)) vasim_50_ste_252 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_251 }),
                .match(vasim_50_w_match_252) ,
                .active_state(vasim_50_w_out_252));




/*wire vasim_50_w_out_253;
*/

wire vasim_50_lut_match_253;
wire vasim_50_w_match_253;

    
    
    

LUT_Match_vasim_50_253 #(8) lut_match_vasim_50_253(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_253));


assign vasim_50_w_match_253 = vasim_50_lut_match_253 ;

STE #(.fan_in(1)) vasim_50_ste_253 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_252 }),
                .match(vasim_50_w_match_253) ,
                .active_state(vasim_50_w_out_253));




/*wire vasim_50_w_out_254;
*/

wire vasim_50_lut_match_254;
wire vasim_50_w_match_254;

    
    
    

LUT_Match_vasim_50_254 #(8) lut_match_vasim_50_254(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_254));


assign vasim_50_w_match_254 = vasim_50_lut_match_254 ;

STE #(.fan_in(1)) vasim_50_ste_254 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_253 }),
                .match(vasim_50_w_match_254) ,
                .active_state(vasim_50_w_out_254));




/*wire vasim_50_w_out_255;
*/

wire vasim_50_lut_match_255;
wire vasim_50_w_match_255;

    
    
    

LUT_Match_vasim_50_255 #(8) lut_match_vasim_50_255(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_255));


assign vasim_50_w_match_255 = vasim_50_lut_match_255 ;

STE #(.fan_in(1)) vasim_50_ste_255 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_254 }),
                .match(vasim_50_w_match_255) ,
                .active_state(vasim_50_w_out_255));




/*wire vasim_50_w_out_256;
*/

wire vasim_50_lut_match_256;
wire vasim_50_w_match_256;

    
    
    

LUT_Match_vasim_50_256 #(8) lut_match_vasim_50_256(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_256));


assign vasim_50_w_match_256 = vasim_50_lut_match_256 ;

STE #(.fan_in(1)) vasim_50_ste_256 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_255 }),
                .match(vasim_50_w_match_256) ,
                .active_state(vasim_50_w_out_256));




/*wire vasim_50_w_out_257;
*/

wire vasim_50_lut_match_257;
wire vasim_50_w_match_257;

    
    
    

LUT_Match_vasim_50_257 #(8) lut_match_vasim_50_257(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_257));


assign vasim_50_w_match_257 = vasim_50_lut_match_257 ;

STE #(.fan_in(1)) vasim_50_ste_257 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_256 }),
                .match(vasim_50_w_match_257) ,
                .active_state(vasim_50_w_out_257));




/*wire vasim_50_w_out_258;
*/

wire vasim_50_lut_match_258;
wire vasim_50_w_match_258;

    
    
    

LUT_Match_vasim_50_258 #(8) lut_match_vasim_50_258(
                .clk(clk),
                .symbols(symbols),
                .match(vasim_50_lut_match_258));


assign vasim_50_w_match_258 = vasim_50_lut_match_258 ;

STE #(.fan_in(1)) vasim_50_ste_258 (
                .clk(clk),
                .run(run),
                .reset(reset),
                .income_edges({ vasim_50_w_out_257 }),
                .match(vasim_50_w_match_258) ,
                .active_state(vasim_50_w_out_258));




endmodule

